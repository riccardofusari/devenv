
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_REGISTER_FILE_WINDOWING is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_REGISTER_FILE_WINDOWING;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_REGISTER_FILE_WINDOWING.all;

entity REGISTER_FILE_WINDOWING_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end REGISTER_FILE_WINDOWING_DW01_add_0;

architecture SYN_cla of REGISTER_FILE_WINDOWING_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244 : std_logic;

begin
   
   U2 : OR2_X1 port map( A1 => B(15), A2 => A(15), ZN => n194);
   U3 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n12);
   U4 : AND2_X1 port map( A1 => n36, A2 => n104, ZN => n96);
   U5 : OR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n159);
   U6 : OR2_X1 port map( A1 => B(17), A2 => A(17), ZN => n158);
   U7 : INV_X1 port map( A => n12, ZN => n226);
   U8 : INV_X1 port map( A => n11, ZN => n80);
   U9 : AND2_X1 port map( A1 => n80, A2 => n79, ZN => n1);
   U10 : AND3_X1 port map( A1 => n113, A2 => n111, A3 => n118, ZN => n2);
   U11 : NOR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n3);
   U12 : AND2_X1 port map( A1 => n110, A2 => n109, ZN => n4);
   U13 : NAND2_X1 port map( A1 => n153, A2 => n7, ZN => n5);
   U14 : AND2_X1 port map( A1 => n5, A2 => n6, ZN => n150);
   U15 : OR2_X1 port map( A1 => n139, A2 => n140, ZN => n6);
   U16 : AND2_X1 port map( A1 => n154, A2 => n143, ZN => n7);
   U17 : OR2_X1 port map( A1 => n161, A2 => n31, ZN => n157);
   U18 : CLKBUF_X1 port map( A => n237, Z => n8);
   U19 : CLKBUF_X1 port map( A => n62, Z => n9);
   U20 : NAND2_X1 port map( A1 => n119, A2 => n2, ZN => n108);
   U21 : NAND2_X1 port map( A1 => n108, A2 => n4, ZN => n105);
   U22 : OR2_X1 port map( A1 => B(27), A2 => A(27), ZN => n113);
   U23 : OR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n62);
   U24 : CLKBUF_X1 port map( A => n206, Z => n10);
   U25 : CLKBUF_X1 port map( A => n69, Z => n16);
   U26 : NOR2_X1 port map( A1 => B(5), A2 => A(5), ZN => n11);
   U27 : NOR2_X1 port map( A1 => B(5), A2 => A(5), ZN => n17);
   U28 : INV_X1 port map( A => n18, ZN => n68);
   U29 : CLKBUF_X1 port map( A => B(7), Z => n13);
   U30 : CLKBUF_X1 port map( A => n221, Z => n14);
   U31 : AND3_X1 port map( A1 => n138, A2 => n136, A3 => n143, ZN => n15);
   U32 : OR2_X1 port map( A1 => B(6), A2 => A(6), ZN => n69);
   U33 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n18);
   U34 : OR2_X2 port map( A1 => B(19), A2 => A(19), ZN => n160);
   U35 : OR2_X2 port map( A1 => B(4), A2 => A(4), ZN => n79);
   U36 : OR2_X1 port map( A1 => n13, A2 => A(7), ZN => n19);
   U37 : XNOR2_X1 port map( A => n40, B => n20, ZN => SUM(10));
   U38 : NAND2_X1 port map( A1 => n226, A2 => n14, ZN => n20);
   U39 : XNOR2_X1 port map( A => n70, B => n21, ZN => SUM(6));
   U40 : NAND2_X1 port map( A1 => n16, A2 => n68, ZN => n21);
   U41 : OR2_X2 port map( A1 => B(23), A2 => A(23), ZN => n138);
   U42 : INV_X1 port map( A => n217, ZN => n22);
   U43 : AND2_X1 port map( A1 => n220, A2 => n219, ZN => n35);
   U44 : XNOR2_X1 port map( A => n213, B => n23, ZN => SUM(14));
   U45 : NAND2_X1 port map( A1 => n192, A2 => n195, ZN => n23);
   U46 : XNOR2_X1 port map( A => n24, B => n25, ZN => SUM(7));
   U47 : AND2_X1 port map( A1 => n67, A2 => n68, ZN => n24);
   U48 : AND2_X1 port map( A1 => n19, A2 => n72, ZN => n25);
   U49 : OAI21_X1 port map( B1 => n22, B2 => n216, A => n198, ZN => n26);
   U50 : OAI21_X1 port map( B1 => n35, B2 => n216, A => n198, ZN => n215);
   U51 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => n27);
   U52 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => n133);
   U53 : AND2_X1 port map( A1 => n15, A2 => n154, ZN => n28);
   U54 : XNOR2_X1 port map( A => n96, B => n29, ZN => SUM(29));
   U55 : AND2_X1 port map( A1 => n97, A2 => n98, ZN => n29);
   U56 : OR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n30);
   U57 : NAND3_X1 port map( A1 => n160, A2 => n159, A3 => n158, ZN => n31);
   U58 : NAND2_X1 port map( A1 => n130, A2 => n34, ZN => n32);
   U59 : AND2_X1 port map( A1 => n32, A2 => n33, ZN => n128);
   U60 : OR2_X1 port map( A1 => n114, A2 => n115, ZN => n33);
   U61 : AND2_X1 port map( A1 => n131, A2 => n118, ZN => n34);
   U62 : OR2_X1 port map( A1 => B(13), A2 => A(13), ZN => n203);
   U63 : NAND2_X1 port map( A1 => n105, A2 => n106, ZN => n36);
   U64 : CLKBUF_X1 port map( A => n227, Z => n37);
   U65 : XNOR2_X1 port map( A => n38, B => n237, ZN => SUM(4));
   U66 : AND2_X1 port map( A1 => n78, A2 => n79, ZN => n38);
   U67 : AND2_X1 port map( A1 => n222, A2 => n48, ZN => n39);
   U68 : OAI21_X1 port map( B1 => n37, B2 => n46, A => n63, ZN => n40);
   U69 : OAI21_X1 port map( B1 => n8, B2 => n209, A => n206, ZN => n41);
   U70 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n42);
   U71 : NAND3_X1 port map( A1 => n133, A2 => n134, A3 => n135, ZN => n43);
   U72 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n44);
   U73 : OR2_X1 port map( A1 => n186, A2 => n187, ZN => n45);
   U74 : NAND2_X1 port map( A1 => n188, A2 => n45, ZN => n183);
   U75 : AND2_X1 port map( A1 => n233, A2 => n65, ZN => n46);
   U76 : OR2_X1 port map( A1 => n210, A2 => n211, ZN => n50);
   U77 : INV_X1 port map( A => n8, ZN => n47);
   U78 : AND3_X1 port map( A1 => n221, A2 => n9, A3 => n66, ZN => n48);
   U79 : AND2_X1 port map( A1 => n222, A2 => n48, ZN => n54);
   U80 : NAND2_X1 port map( A1 => n210, A2 => n211, ZN => n49);
   U81 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => SUM(15));
   U82 : NAND3_X1 port map( A1 => n71, A2 => n16, A3 => n1, ZN => n209);
   U83 : XOR2_X1 port map( A => n51, B => n149, Z => SUM(22));
   U84 : AND2_X1 port map( A1 => n136, A2 => n142, ZN => n51);
   U85 : XOR2_X1 port map( A => n52, B => n129, Z => SUM(25));
   U86 : AND2_X1 port map( A1 => n118, A2 => n116, ZN => n52);
   U87 : OR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n221);
   U88 : AND2_X1 port map( A1 => n173, A2 => n238, ZN => SUM(0));
   U89 : OR2_X1 port map( A1 => B(22), A2 => A(22), ZN => n136);
   U90 : OR2_X1 port map( A1 => B(21), A2 => A(21), ZN => n143);
   U91 : OR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n118);
   U92 : OR2_X1 port map( A1 => B(26), A2 => A(26), ZN => n111);
   U93 : OR2_X1 port map( A1 => B(29), A2 => A(29), ZN => n98);
   U94 : INV_X1 port map( A => B(0), ZN => n243);
   U95 : XNOR2_X1 port map( A => n105, B => n107, ZN => SUM(28));
   U96 : OAI21_X1 port map( B1 => n8, B2 => n209, A => n206, ZN => n64);
   U97 : OAI21_X1 port map( B1 => n46, B2 => n37, A => n63, ZN => n232);
   U98 : OAI21_X1 port map( B1 => n3, B2 => n173, A => n101, ZN => n241);
   U99 : OAI21_X1 port map( B1 => n73, B2 => n11, A => n74, ZN => n70);
   U100 : OAI21_X1 port map( B1 => n223, B2 => n42, A => n224, ZN => n205);
   U101 : AOI21_X1 port map( B1 => n225, B2 => n221, A => n12, ZN => n223);
   U102 : OAI21_X1 port map( B1 => n227, B2 => n65, A => n63, ZN => n225);
   U103 : XNOR2_X1 port map( A => n99, B => n86, ZN => SUM(2));
   U104 : NAND2_X1 port map( A1 => n103, A2 => n85, ZN => n99);
   U105 : AOI21_X1 port map( B1 => n39, B2 => n204, A => n205, ZN => n186);
   U106 : NOR2_X1 port map( A1 => n190, A2 => n189, ZN => n188);
   U107 : NAND2_X1 port map( A1 => n161, A2 => n169, ZN => n181);
   U108 : NAND2_X1 port map( A1 => n180, A2 => n170, ZN => n178);
   U109 : NAND2_X1 port map( A1 => n158, A2 => n181, ZN => n180);
   U110 : XNOR2_X1 port map( A => n179, B => n178, ZN => SUM(18));
   U111 : NAND2_X1 port map( A1 => n165, A2 => n159, ZN => n179);
   U112 : NAND2_X1 port map( A1 => n195, A2 => n196, ZN => n191);
   U113 : OAI21_X1 port map( B1 => n197, B2 => n198, A => n199, ZN => n196);
   U114 : XOR2_X1 port map( A => n41, B => n55, Z => SUM(8));
   U115 : AND2_X1 port map( A1 => n65, A2 => n66, ZN => n55);
   U116 : XOR2_X1 port map( A => n56, B => n26, Z => SUM(13));
   U117 : AND2_X1 port map( A1 => n199, A2 => n203, ZN => n56);
   U118 : INV_X1 port map( A => n173, ZN => n102);
   U119 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => n86);
   U120 : NAND2_X1 port map( A1 => n30, A2 => n102, ZN => n100);
   U121 : NAND2_X1 port map( A1 => n171, A2 => n160, ZN => n174);
   U122 : NAND2_X1 port map( A1 => n80, A2 => n74, ZN => n76);
   U123 : NAND2_X1 port map( A1 => n9, A2 => n63, ZN => n60);
   U124 : NOR2_X1 port map( A1 => n162, A2 => n163, ZN => n156);
   U125 : NAND2_X1 port map( A1 => n150, A2 => n141, ZN => n149);
   U126 : NAND2_X1 port map( A1 => n144, A2 => n140, ZN => n151);
   U127 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n91);
   U128 : OAI211_X1 port map( C1 => n139, C2 => n140, A => n141, B => n142, ZN 
                           => n137);
   U129 : OAI211_X1 port map( C1 => n114, C2 => n115, A => n116, B => n117, ZN 
                           => n112);
   U130 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n81);
   U131 : NAND2_X1 port map( A1 => n128, A2 => n116, ZN => n125);
   U132 : NAND2_X1 port map( A1 => n120, A2 => n115, ZN => n129);
   U133 : XNOR2_X1 port map( A => n125, B => n127, ZN => SUM(26));
   U134 : NAND2_X1 port map( A1 => n111, A2 => n117, ZN => n127);
   U135 : NAND2_X1 port map( A1 => n134, A2 => n138, ZN => n145);
   U136 : OAI21_X1 port map( B1 => n147, B2 => n148, A => n142, ZN => n146);
   U137 : NAND2_X1 port map( A1 => n198, A2 => n202, ZN => n218);
   U138 : XNOR2_X1 port map( A => n121, B => n122, ZN => SUM(27));
   U139 : NOR2_X1 port map( A1 => n123, A2 => n124, ZN => n122);
   U140 : AOI21_X1 port map( B1 => n125, B2 => n111, A => n126, ZN => n121);
   U141 : XOR2_X1 port map( A => n89, B => n90, Z => SUM(31));
   U142 : XNOR2_X1 port map( A => n182, B => n181, ZN => SUM(17));
   U143 : NAND2_X1 port map( A1 => n170, A2 => n158, ZN => n182);
   U144 : AOI21_X1 port map( B1 => n164, B2 => n165, A => n166, ZN => n163);
   U145 : NAND2_X1 port map( A1 => n159, A2 => n167, ZN => n164);
   U146 : OAI21_X1 port map( B1 => n168, B2 => n169, A => n170, ZN => n167);
   U147 : NAND2_X1 port map( A1 => n169, A2 => n184, ZN => n185);
   U148 : NAND2_X1 port map( A1 => n143, A2 => n141, ZN => n152);
   U149 : NAND2_X1 port map( A1 => n154, A2 => n140, ZN => n155);
   U150 : XNOR2_X1 port map( A => n172, B => n102, ZN => SUM(1));
   U151 : NAND2_X1 port map( A1 => n30, A2 => n101, ZN => n172);
   U152 : NAND2_X1 port map( A1 => n10, A2 => n207, ZN => n204);
   U153 : NAND2_X1 port map( A1 => n131, A2 => n115, ZN => n132);
   U154 : NAND2_X1 port map( A1 => n104, A2 => n106, ZN => n107);
   U155 : OR2_X1 port map( A1 => B(3), A2 => A(3), ZN => n87);
   U156 : OR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n222);
   U157 : OR2_X1 port map( A1 => B(2), A2 => A(2), ZN => n103);
   U158 : NAND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n173);
   U159 : OR2_X2 port map( A1 => B(14), A2 => A(14), ZN => n195);
   U160 : XNOR2_X1 port map( A => n91, B => n93, ZN => SUM(30));
   U161 : NAND2_X1 port map( A1 => n92, A2 => n94, ZN => n93);
   U162 : NAND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n94);
   U163 : NAND2_X1 port map( A1 => B(13), A2 => A(13), ZN => n199);
   U164 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n63);
   U165 : NAND2_X1 port map( A1 => n243, A2 => n244, ZN => n238);
   U166 : INV_X1 port map( A => A(0), ZN => n244);
   U167 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n192);
   U168 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n65);
   U169 : NAND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n198);
   U170 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n66);
   U171 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n171);
   U172 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n165);
   U173 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n170);
   U174 : OR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n202);
   U175 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n142);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => A(26), ZN => n117);
   U177 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n169);
   U178 : NAND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n134);
   U179 : OR2_X1 port map( A1 => B(16), A2 => A(16), ZN => n184);
   U180 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n141);
   U181 : NAND2_X1 port map( A1 => B(27), A2 => A(27), ZN => n109);
   U182 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n116);
   U183 : OR2_X1 port map( A1 => B(20), A2 => A(20), ZN => n154);
   U184 : OR2_X1 port map( A1 => B(30), A2 => A(30), ZN => n92);
   U185 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n140);
   U186 : OR2_X1 port map( A1 => B(24), A2 => A(24), ZN => n131);
   U187 : NAND2_X1 port map( A1 => B(24), A2 => A(24), ZN => n115);
   U188 : OR2_X1 port map( A1 => B(28), A2 => A(28), ZN => n106);
   U189 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n97);
   U190 : NAND2_X1 port map( A1 => B(28), A2 => A(28), ZN => n104);
   U191 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n90);
   U192 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => n57);
   U193 : OAI21_X1 port map( B1 => n239, B2 => n240, A => n88, ZN => n208);
   U194 : OAI21_X1 port map( B1 => n77, B2 => n237, A => n78, ZN => n75);
   U195 : NAND2_X1 port map( A1 => B(4), A2 => A(4), ZN => n78);
   U196 : XNOR2_X1 port map( A => n152, B => n151, ZN => SUM(21));
   U197 : XNOR2_X1 port map( A => n155, B => n153, ZN => SUM(20));
   U198 : NAND2_X1 port map( A1 => n153, A2 => n154, ZN => n144);
   U199 : NAND2_X1 port map( A1 => n200, A2 => n194, ZN => n210);
   U200 : NAND4_X1 port map( A1 => n194, A2 => n203, A3 => n195, A4 => n202, ZN
                           => n187);
   U201 : AOI21_X1 port map( B1 => n191, B2 => n192, A => n193, ZN => n190);
   U202 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => n74);
   U203 : OAI21_X1 port map( B1 => n214, B2 => n197, A => n199, ZN => n58);
   U204 : OAI21_X1 port map( B1 => n214, B2 => n197, A => n199, ZN => n213);
   U205 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n85);
   U206 : XNOR2_X1 port map( A => n43, B => n132, ZN => SUM(24));
   U207 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n120);
   U208 : NAND2_X1 port map( A1 => n156, A2 => n157, ZN => n153);
   U209 : NAND2_X1 port map( A1 => n183, A2 => n184, ZN => n161);
   U210 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n200);
   U211 : NOR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n59);
   U212 : AOI21_X1 port map( B1 => n69, B2 => n236, A => n18, ZN => n235);
   U213 : OAI21_X1 port map( B1 => n17, B2 => n78, A => n74, ZN => n236);
   U214 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n71);
   U215 : NAND2_X1 port map( A1 => n212, A2 => n192, ZN => n211);
   U216 : NAND2_X1 port map( A1 => n58, A2 => n195, ZN => n212);
   U217 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => n88);
   U218 : XNOR2_X1 port map( A => n217, B => n218, ZN => SUM(12));
   U219 : NAND2_X1 port map( A1 => n220, A2 => n219, ZN => n217);
   U220 : XNOR2_X1 port map( A => n60, B => n61, ZN => SUM(9));
   U221 : NAND2_X1 port map( A1 => n233, A2 => n65, ZN => n61);
   U222 : OAI21_X1 port map( B1 => n59, B2 => n235, A => n72, ZN => n234);
   U223 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n101);
   U224 : AOI21_X1 port map( B1 => n241, B2 => n103, A => n242, ZN => n239);
   U225 : NAND2_X1 port map( A1 => n224, A2 => n222, ZN => n228);
   U226 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n224);
   U227 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n72);
   U228 : NAND2_X1 port map( A1 => n16, A2 => n70, ZN => n67);
   U229 : XNOR2_X1 port map( A => n75, B => n76, ZN => SUM(5));
   U230 : NAND2_X1 port map( A1 => n64, A2 => n66, ZN => n233);
   U231 : NAND2_X1 port map( A1 => n54, A2 => n41, ZN => n220);
   U232 : NAND2_X1 port map( A1 => n201, A2 => n47, ZN => n207);
   U233 : INV_X1 port map( A => n75, ZN => n73);
   U234 : INV_X1 port map( A => n79, ZN => n77);
   U235 : XNOR2_X1 port map( A => n81, B => n82, ZN => SUM(3));
   U236 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U237 : INV_X1 port map( A => n86, ZN => n83);
   U238 : AOI21_X1 port map( B1 => n44, B2 => n92, A => n57, ZN => n89);
   U239 : INV_X1 port map( A => n98, ZN => n95);
   U240 : NAND3_X1 port map( A1 => n111, A2 => n112, A3 => n113, ZN => n110);
   U241 : INV_X1 port map( A => n118, ZN => n114);
   U242 : INV_X1 port map( A => n120, ZN => n119);
   U243 : INV_X1 port map( A => n109, ZN => n124);
   U244 : INV_X1 port map( A => n113, ZN => n123);
   U245 : INV_X1 port map( A => n117, ZN => n126);
   U246 : NAND3_X1 port map( A1 => n133, A2 => n134, A3 => n135, ZN => n130);
   U247 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n138, ZN => n135);
   U248 : INV_X1 port map( A => n143, ZN => n139);
   U249 : XNOR2_X1 port map( A => n145, B => n146, ZN => SUM(23));
   U250 : INV_X1 port map( A => n136, ZN => n148);
   U251 : INV_X1 port map( A => n149, ZN => n147);
   U252 : INV_X1 port map( A => n160, ZN => n166);
   U253 : INV_X1 port map( A => n158, ZN => n168);
   U254 : INV_X1 port map( A => n171, ZN => n162);
   U255 : XNOR2_X1 port map( A => n175, B => n174, ZN => SUM(19));
   U256 : OAI21_X1 port map( B1 => n176, B2 => n177, A => n165, ZN => n175);
   U257 : INV_X1 port map( A => n159, ZN => n177);
   U258 : INV_X1 port map( A => n178, ZN => n176);
   U259 : XNOR2_X1 port map( A => n185, B => n183, ZN => SUM(16));
   U260 : INV_X1 port map( A => n194, ZN => n193);
   U261 : INV_X1 port map( A => n200, ZN => n189);
   U262 : INV_X1 port map( A => n209, ZN => n201);
   U263 : INV_X1 port map( A => n203, ZN => n197);
   U264 : INV_X1 port map( A => n215, ZN => n214);
   U265 : INV_X1 port map( A => n202, ZN => n216);
   U266 : INV_X1 port map( A => n205, ZN => n219);
   U267 : XNOR2_X1 port map( A => n229, B => n228, ZN => SUM(11));
   U268 : OAI21_X1 port map( B1 => n230, B2 => n231, A => n226, ZN => n229);
   U269 : INV_X1 port map( A => n14, ZN => n231);
   U270 : INV_X1 port map( A => n232, ZN => n230);
   U271 : INV_X1 port map( A => n234, ZN => n206);
   U272 : INV_X1 port map( A => n103, ZN => n84);
   U273 : INV_X1 port map( A => n208, ZN => n237);
   U274 : INV_X1 port map( A => n87, ZN => n240);
   U275 : INV_X1 port map( A => n85, ZN => n242);
   U276 : INV_X1 port map( A => n62, ZN => n227);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_REGISTER_FILE_WINDOWING.all;

entity REGISTER_FILE_WINDOWING_DW01_addsub_2 is

   port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (31 downto 0);  CO : out std_logic);

end REGISTER_FILE_WINDOWING_DW01_addsub_2;

architecture SYN_cla of REGISTER_FILE_WINDOWING_DW01_addsub_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261 : std_logic;

begin
   
   U2 : INV_X1 port map( A => n13, ZN => n219);
   U3 : BUF_X2 port map( A => n78, Z => n40);
   U4 : AND2_X1 port map( A1 => n130, A2 => n136, ZN => n1);
   U5 : AND2_X1 port map( A1 => n103, A2 => n110, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n11, B2 => n208, A => n238, ZN => n3);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n208, A => n238, ZN => n47);
   U8 : XNOR2_X1 port map( A => n9, B => n4, ZN => SUM(13));
   U9 : NAND2_X1 port map( A1 => n187, A2 => n201, ZN => n4);
   U10 : CLKBUF_X1 port map( A => n206, Z => n19);
   U11 : XNOR2_X1 port map( A => n67, B => n18, ZN => SUM(4));
   U12 : CLKBUF_X1 port map( A => n202, Z => n5);
   U13 : CLKBUF_X1 port map( A => A(0), Z => n6);
   U14 : OR2_X1 port map( A1 => n206, A2 => n29, ZN => n18);
   U15 : INV_X1 port map( A => n40, ZN => n38);
   U16 : AND2_X1 port map( A1 => n90, A2 => n14, ZN => n7);
   U17 : BUF_X1 port map( A => n10, Z => n14);
   U18 : INV_X2 port map( A => n40, ZN => n39);
   U19 : CLKBUF_X1 port map( A => n71, Z => n8);
   U20 : OAI21_X1 port map( B1 => n13, B2 => n218, A => n188, ZN => n9);
   U21 : NAND2_X1 port map( A1 => n165, A2 => A(1), ZN => n10);
   U22 : NOR2_X1 port map( A1 => n206, A2 => n29, ZN => n11);
   U23 : AND2_X1 port map( A1 => n64, A2 => n65, ZN => n12);
   U24 : AND2_X2 port map( A1 => n31, A2 => n222, ZN => n13);
   U25 : AND2_X1 port map( A1 => n243, A2 => n92, ZN => n15);
   U26 : AND2_X1 port map( A1 => n244, A2 => n15, ZN => n29);
   U27 : AND2_X1 port map( A1 => n253, A2 => n255, ZN => n16);
   U28 : OR2_X1 port map( A1 => n29, A2 => n206, ZN => n17);
   U29 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => n20);
   U30 : NAND2_X1 port map( A1 => n247, A2 => n250, ZN => n21);
   U31 : AND2_X1 port map( A1 => n216, A2 => n187, ZN => n22);
   U32 : AND2_X1 port map( A1 => n20, A2 => n49, ZN => n23);
   U33 : XNOR2_X1 port map( A => n89, B => n73, ZN => SUM(2));
   U34 : OAI21_X1 port map( B1 => n13, B2 => n218, A => n188, ZN => n24);
   U35 : AND2_X1 port map( A1 => n236, A2 => n49, ZN => n25);
   U36 : CLKBUF_X1 port map( A => n41, Z => n36);
   U37 : NOR2_X1 port map( A1 => n26, A2 => n27, ZN => n97);
   U38 : NOR2_X1 port map( A1 => n107, A2 => n108, ZN => n26);
   U39 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN 
                           => n27);
   U40 : XOR2_X1 port map( A => n28, B => n144, Z => SUM(21));
   U41 : AND2_X1 port map( A1 => n132, A2 => n135, ZN => n28);
   U42 : BUF_X1 port map( A => n36, Z => n35);
   U43 : BUF_X1 port map( A => n36, Z => n34);
   U44 : OAI21_X1 port map( B1 => n181, B2 => n182, A => n183, ZN => n178);
   U45 : INV_X1 port map( A => n203, ZN => n181);
   U46 : OAI21_X1 port map( B1 => n204, B2 => n205, A => n31, ZN => n203);
   U47 : NOR2_X1 port map( A1 => n193, A2 => n194, ZN => n184);
   U48 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n50);
   U49 : OAI21_X1 port map( B1 => n12, B2 => n59, A => n60, ZN => n55);
   U50 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => n58);
   U51 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => n68);
   U52 : NAND2_X1 port map( A1 => n61, A2 => n60, ZN => n63);
   U53 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => n89);
   U54 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => n228);
   U55 : XNOR2_X1 port map( A => n37, B => n234, ZN => SUM(10));
   U56 : NAND2_X1 port map( A1 => n226, A2 => n223, ZN => n234);
   U57 : NAND2_X1 port map( A1 => n190, A2 => n199, ZN => n210);
   U58 : INV_X1 port map( A => ADD_SUB, ZN => n78);
   U59 : XNOR2_X1 port map( A => n40, B => n30, ZN => SUM(0));
   U60 : AND2_X1 port map( A1 => n192, A2 => n164, ZN => n30);
   U61 : AND2_X1 port map( A1 => n72, A2 => n74, ZN => n244);
   U62 : XNOR2_X1 port map( A => n215, B => n213, ZN => SUM(14));
   U63 : NAND2_X1 port map( A1 => n189, A2 => n200, ZN => n215);
   U64 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n42);
   U65 : INV_X1 port map( A => ADD_SUB, ZN => n261);
   U66 : NAND4_X1 port map( A1 => n223, A2 => n224, A3 => n44, A4 => n48, ZN =>
                           n205);
   U67 : NAND4_X1 port map( A1 => n66, A2 => n61, A3 => n54, A4 => n56, ZN => 
                           n208);
   U68 : AND4_X1 port map( A1 => n225, A2 => n45, A3 => n49, A4 => n226, ZN => 
                           n31);
   U69 : NAND2_X1 port map( A1 => n155, A2 => n161, ZN => n166);
   U70 : NAND2_X1 port map( A1 => n150, A2 => n158, ZN => n174);
   U71 : NAND2_X1 port map( A1 => n173, A2 => n157, ZN => n170);
   U72 : NAND2_X1 port map( A1 => n160, A2 => n174, ZN => n173);
   U73 : NAND2_X1 port map( A1 => n177, A2 => n178, ZN => n150);
   U74 : NAND4_X1 port map( A1 => n199, A2 => n200, A3 => n201, A4 => n202, ZN 
                           => n182);
   U75 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => n46);
   U76 : XNOR2_X1 port map( A => n221, B => n219, ZN => SUM(12));
   U77 : NAND2_X1 port map( A1 => n188, A2 => n5, ZN => n221);
   U78 : XNOR2_X1 port map( A => n172, B => n170, ZN => SUM(18));
   U79 : NAND2_X1 port map( A1 => n156, A2 => n159, ZN => n172);
   U80 : XNOR2_X1 port map( A => n176, B => n174, ZN => SUM(17));
   U81 : NAND2_X1 port map( A1 => n157, A2 => n160, ZN => n176);
   U82 : NAND4_X1 port map( A1 => n187, A2 => n188, A3 => n189, A4 => n190, ZN 
                           => n186);
   U83 : OAI21_X1 port map( B1 => n150, B2 => n151, A => n152, ZN => n146);
   U84 : NOR2_X1 port map( A1 => n153, A2 => n154, ZN => n152);
   U85 : NAND2_X1 port map( A1 => n157, A2 => n158, ZN => n153);
   U86 : XNOR2_X1 port map( A => n137, B => n1, ZN => SUM(23));
   U87 : AOI21_X1 port map( B1 => n134, B2 => n139, A => n140, ZN => n137);
   U88 : NAND2_X1 port map( A1 => n125, A2 => n133, ZN => n144);
   U89 : NAND2_X1 port map( A1 => n143, A2 => n132, ZN => n139);
   U90 : NAND2_X1 port map( A1 => n135, A2 => n144, ZN => n143);
   U91 : NAND2_X1 port map( A1 => n145, A2 => n146, ZN => n125);
   U92 : XNOR2_X1 port map( A => n139, B => n141, ZN => SUM(22));
   U93 : NAND2_X1 port map( A1 => n134, A2 => n131, ZN => n141);
   U94 : OAI21_X1 port map( B1 => n125, B2 => n126, A => n127, ZN => n121);
   U95 : NOR2_X1 port map( A1 => n128, A2 => n129, ZN => n127);
   U96 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => n128);
   U97 : XNOR2_X1 port map( A => n112, B => n2, ZN => SUM(27));
   U98 : AOI21_X1 port map( B1 => n111, B2 => n114, A => n115, ZN => n112);
   U99 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => n119);
   U100 : NAND2_X1 port map( A1 => n118, A2 => n105, ZN => n114);
   U101 : NAND2_X1 port map( A1 => n109, A2 => n119, ZN => n118);
   U102 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => n107);
   U103 : XNOR2_X1 port map( A => n114, B => n116, ZN => SUM(26));
   U104 : NAND2_X1 port map( A1 => n111, A2 => n104, ZN => n116);
   U105 : NAND2_X1 port map( A1 => n158, A2 => n177, ZN => n180);
   U106 : XOR2_X1 port map( A => n32, B => n119, Z => SUM(25));
   U107 : AND2_X1 port map( A1 => n105, A2 => n109, ZN => n32);
   U108 : XNOR2_X1 port map( A => n146, B => n148, ZN => SUM(20));
   U109 : NAND2_X1 port map( A1 => n145, A2 => n133, ZN => n148);
   U110 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n80);
   U111 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n96);
   U112 : XNOR2_X1 port map( A => n80, B => n83, ZN => SUM(30));
   U113 : NAND2_X1 port map( A1 => n82, A2 => n79, ZN => n83);
   U114 : XNOR2_X1 port map( A => n121, B => n123, ZN => SUM(24));
   U115 : NAND2_X1 port map( A1 => n120, A2 => n106, ZN => n123);
   U116 : XOR2_X1 port map( A => n85, B => n94, Z => SUM(29));
   U117 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n94);
   U118 : NAND2_X1 port map( A1 => n155, A2 => n156, ZN => n154);
   U119 : XOR2_X1 port map( A => n97, B => n101, Z => SUM(28));
   U120 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n101);
   U121 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n129);
   U122 : NAND2_X1 port map( A1 => A(6), A2 => n38, ZN => n53);
   U123 : NAND2_X1 port map( A1 => A(4), A2 => n38, ZN => n65);
   U124 : NAND2_X1 port map( A1 => A(5), A2 => n38, ZN => n60);
   U125 : NAND2_X1 port map( A1 => A(7), A2 => n38, ZN => n57);
   U126 : NAND2_X1 port map( A1 => n78, A2 => n237, ZN => n48);
   U127 : INV_X1 port map( A => A(8), ZN => n237);
   U128 : NAND2_X1 port map( A1 => n247, A2 => n250, ZN => n74);
   U129 : INV_X1 port map( A => A(3), ZN => n250);
   U130 : NAND2_X1 port map( A1 => n78, A2 => n256, ZN => n44);
   U131 : INV_X1 port map( A => A(9), ZN => n256);
   U132 : NAND2_X1 port map( A1 => n78, A2 => n233, ZN => n224);
   U133 : INV_X1 port map( A => A(11), ZN => n233);
   U134 : NAND2_X1 port map( A1 => n78, A2 => n257, ZN => n223);
   U135 : INV_X1 port map( A => A(10), ZN => n257);
   U136 : INV_X1 port map( A => A(7), ZN => n239);
   U137 : INV_X1 port map( A => A(5), ZN => n241);
   U138 : INV_X1 port map( A => A(6), ZN => n240);
   U139 : NAND2_X1 port map( A1 => A(9), A2 => n39, ZN => n45);
   U140 : NAND2_X1 port map( A1 => A(8), A2 => n39, ZN => n49);
   U141 : INV_X1 port map( A => A(4), ZN => n242);
   U142 : NAND2_X1 port map( A1 => A(10), A2 => n39, ZN => n226);
   U143 : NAND2_X1 port map( A1 => A(3), A2 => n246, ZN => n75);
   U144 : NAND2_X1 port map( A1 => A(11), A2 => n39, ZN => n225);
   U145 : NAND2_X1 port map( A1 => n41, A2 => n227, ZN => n202);
   U146 : INV_X1 port map( A => A(12), ZN => n227);
   U147 : NAND2_X1 port map( A1 => n41, A2 => n220, ZN => n201);
   U148 : INV_X1 port map( A => A(13), ZN => n220);
   U149 : NAND2_X1 port map( A1 => n40, A2 => n217, ZN => n200);
   U150 : INV_X1 port map( A => A(14), ZN => n217);
   U151 : NAND2_X1 port map( A1 => n40, A2 => n214, ZN => n199);
   U152 : INV_X1 port map( A => A(15), ZN => n214);
   U153 : NAND2_X1 port map( A1 => A(12), A2 => n39, ZN => n188);
   U154 : NAND2_X1 port map( A1 => A(15), A2 => n39, ZN => n190);
   U155 : NAND2_X1 port map( A1 => A(13), A2 => n198, ZN => n187);
   U156 : NAND2_X1 port map( A1 => A(14), A2 => n198, ZN => n189);
   U157 : NAND2_X1 port map( A1 => n36, A2 => n209, ZN => n177);
   U158 : INV_X1 port map( A => A(16), ZN => n209);
   U159 : NAND2_X1 port map( A1 => A(16), A2 => n39, ZN => n158);
   U160 : NAND2_X1 port map( A1 => A(18), A2 => n198, ZN => n156);
   U161 : NAND2_X1 port map( A1 => n33, A2 => n179, ZN => n160);
   U162 : INV_X1 port map( A => A(17), ZN => n179);
   U163 : NAND2_X1 port map( A1 => A(17), A2 => n39, ZN => n157);
   U164 : NAND2_X1 port map( A1 => n35, A2 => n175, ZN => n159);
   U165 : INV_X1 port map( A => A(18), ZN => n175);
   U166 : NAND2_X1 port map( A1 => n34, A2 => n171, ZN => n161);
   U167 : INV_X1 port map( A => A(19), ZN => n171);
   U168 : NAND2_X1 port map( A1 => A(19), A2 => n39, ZN => n155);
   U169 : NAND2_X1 port map( A1 => n34, A2 => n149, ZN => n145);
   U170 : INV_X1 port map( A => A(20), ZN => n149);
   U171 : NAND2_X1 port map( A1 => A(22), A2 => n39, ZN => n131);
   U172 : NAND2_X1 port map( A1 => A(20), A2 => n39, ZN => n133);
   U173 : NAND2_X1 port map( A1 => A(23), A2 => n39, ZN => n130);
   U174 : NAND2_X1 port map( A1 => A(21), A2 => n198, ZN => n132);
   U175 : NAND2_X1 port map( A1 => n35, A2 => n147, ZN => n135);
   U176 : INV_X1 port map( A => A(21), ZN => n147);
   U177 : NAND2_X1 port map( A1 => n34, A2 => n142, ZN => n134);
   U178 : INV_X1 port map( A => A(22), ZN => n142);
   U179 : NAND2_X1 port map( A1 => n35, A2 => n138, ZN => n136);
   U180 : INV_X1 port map( A => A(23), ZN => n138);
   U181 : NAND2_X1 port map( A1 => n34, A2 => n124, ZN => n120);
   U182 : INV_X1 port map( A => A(24), ZN => n124);
   U183 : NAND2_X1 port map( A1 => A(24), A2 => n38, ZN => n106);
   U184 : NAND2_X1 port map( A1 => n35, A2 => n122, ZN => n109);
   U185 : INV_X1 port map( A => A(25), ZN => n122);
   U186 : NAND2_X1 port map( A1 => A(25), A2 => n39, ZN => n105);
   U187 : NAND2_X1 port map( A1 => n34, A2 => n113, ZN => n110);
   U188 : INV_X1 port map( A => A(27), ZN => n113);
   U189 : NAND2_X1 port map( A1 => n33, A2 => n117, ZN => n111);
   U190 : INV_X1 port map( A => A(26), ZN => n117);
   U191 : NAND2_X1 port map( A1 => A(26), A2 => n39, ZN => n104);
   U192 : NAND2_X1 port map( A1 => A(27), A2 => n39, ZN => n103);
   U193 : NAND2_X1 port map( A1 => n35, A2 => n102, ZN => n100);
   U194 : INV_X1 port map( A => A(28), ZN => n102);
   U195 : NAND2_X1 port map( A1 => A(28), A2 => n39, ZN => n99);
   U196 : NAND2_X1 port map( A1 => n33, A2 => n95, ZN => n88);
   U197 : INV_X1 port map( A => A(29), ZN => n95);
   U198 : NAND2_X1 port map( A1 => A(29), A2 => n198, ZN => n87);
   U199 : NAND2_X1 port map( A1 => n34, A2 => n84, ZN => n79);
   U200 : INV_X1 port map( A => A(30), ZN => n84);
   U201 : NAND2_X1 port map( A1 => A(30), A2 => n38, ZN => n82);
   U202 : XNOR2_X1 port map( A => n76, B => n77, ZN => SUM(31));
   U203 : NAND2_X1 port map( A1 => n254, A2 => A(2), ZN => n71);
   U204 : INV_X1 port map( A => A(2), ZN => n252);
   U205 : NAND2_X1 port map( A1 => n251, A2 => n252, ZN => n72);
   U206 : XNOR2_X1 port map( A => n69, B => n68, ZN => SUM(3));
   U207 : AOI21_X1 port map( B1 => n197, B2 => n19, A => n207, ZN => n204);
   U208 : BUF_X1 port map( A => n36, Z => n33);
   U209 : XNOR2_X1 port map( A => n93, B => n162, ZN => SUM(1));
   U210 : XNOR2_X1 port map( A => n63, B => n62, ZN => SUM(5));
   U211 : NAND2_X1 port map( A1 => n253, A2 => n255, ZN => n92);
   U212 : NAND2_X1 port map( A1 => n261, A2 => n242, ZN => n66);
   U213 : NAND2_X1 port map( A1 => n261, A2 => n241, ZN => n61);
   U214 : NAND2_X1 port map( A1 => n261, A2 => n240, ZN => n54);
   U215 : NAND2_X1 port map( A1 => n261, A2 => n239, ZN => n56);
   U216 : CLKBUF_X1 port map( A => n78, Z => n41);
   U217 : XNOR2_X1 port map( A => n46, B => n3, ZN => SUM(8));
   U218 : NAND2_X1 port map( A1 => n196, A2 => n47, ZN => n222);
   U219 : NAND2_X1 port map( A1 => n163, A2 => n164, ZN => n93);
   U220 : NAND2_X1 port map( A1 => n198, A2 => n192, ZN => n163);
   U221 : OAI21_X1 port map( B1 => n23, B2 => n235, A => n45, ZN => n37);
   U222 : OAI21_X1 port map( B1 => n25, B2 => n235, A => n45, ZN => n232);
   U223 : NAND2_X1 port map( A1 => n259, A2 => n260, ZN => n192);
   U224 : NAND2_X1 port map( A1 => n216, A2 => n187, ZN => n213);
   U225 : NAND2_X1 port map( A1 => n24, A2 => n201, ZN => n216);
   U226 : NAND2_X1 port map( A1 => n20, A2 => n49, ZN => n43);
   U227 : NAND2_X1 port map( A1 => n6, A2 => n258, ZN => n164);
   U228 : INV_X1 port map( A => A(0), ZN => n260);
   U229 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => n162);
   U230 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => n90);
   U231 : XNOR2_X1 port map( A => n42, B => n43, ZN => SUM(9));
   U232 : XNOR2_X1 port map( A => n51, B => n50, ZN => SUM(7));
   U233 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n51);
   U234 : NAND2_X1 port map( A1 => n17, A2 => n66, ZN => n64);
   U235 : OAI211_X1 port map( C1 => n249, C2 => n248, A => n72, B => n21, ZN =>
                           n245);
   U236 : NAND2_X1 port map( A1 => n90, A2 => n14, ZN => n73);
   U237 : NAND2_X1 port map( A1 => n71, A2 => n10, ZN => n249);
   U238 : NOR2_X1 port map( A1 => n16, A2 => n191, ZN => n185);
   U239 : NOR2_X1 port map( A1 => n16, A2 => n164, ZN => n248);
   U240 : XNOR2_X1 port map( A => n55, B => n58, ZN => SUM(6));
   U241 : NAND2_X1 port map( A1 => n55, A2 => n54, ZN => n52);
   U242 : NAND2_X1 port map( A1 => n165, A2 => A(1), ZN => n91);
   U243 : INV_X1 port map( A => A(1), ZN => n255);
   U244 : NAND2_X1 port map( A1 => n245, A2 => n75, ZN => n206);
   U245 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => n67);
   U246 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n62);
   U247 : NAND4_X1 port map( A1 => n57, A2 => n53, A3 => n60, A4 => n65, ZN => 
                           n207);
   U248 : XNOR2_X1 port map( A => B(3), B => ADD_SUB, ZN => n247);
   U249 : XNOR2_X1 port map( A => B(2), B => ADD_SUB, ZN => n251);
   U250 : XNOR2_X1 port map( A => B(1), B => ADD_SUB, ZN => n253);
   U251 : XNOR2_X1 port map( A => B(0), B => ADD_SUB, ZN => n259);
   U252 : NAND2_X1 port map( A1 => n3, A2 => n48, ZN => n236);
   U253 : INV_X1 port map( A => n61, ZN => n59);
   U254 : OAI21_X1 port map( B1 => n7, B2 => n70, A => n8, ZN => n69);
   U255 : INV_X1 port map( A => n72, ZN => n70);
   U256 : XNOR2_X1 port map( A => A(31), B => n35, ZN => n77);
   U257 : AOI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n76);
   U258 : INV_X1 port map( A => n82, ZN => n81);
   U259 : INV_X1 port map( A => n88, ZN => n86);
   U260 : INV_X1 port map( A => n96, ZN => n85);
   U261 : INV_X1 port map( A => n100, ZN => n98);
   U262 : NAND3_X1 port map( A1 => n109, A2 => n110, A3 => n111, ZN => n108);
   U263 : INV_X1 port map( A => n104, ZN => n115);
   U264 : NAND3_X1 port map( A1 => n134, A2 => n135, A3 => n136, ZN => n126);
   U265 : INV_X1 port map( A => n131, ZN => n140);
   U266 : NAND3_X1 port map( A1 => n159, A2 => n160, A3 => n161, ZN => n151);
   U267 : XNOR2_X1 port map( A => n166, B => n167, ZN => SUM(19));
   U268 : OAI21_X1 port map( B1 => n168, B2 => n169, A => n156, ZN => n167);
   U269 : INV_X1 port map( A => n159, ZN => n169);
   U270 : INV_X1 port map( A => n170, ZN => n168);
   U271 : XNOR2_X1 port map( A => n180, B => n178, ZN => SUM(16));
   U272 : AOI21_X1 port map( B1 => n184, B2 => n185, A => n186, ZN => n183);
   U273 : NAND3_X1 port map( A1 => n192, A2 => n21, A3 => n72, ZN => n191);
   U274 : NAND2_X1 port map( A1 => n195, A2 => n196, ZN => n194);
   U275 : INV_X1 port map( A => n182, ZN => n195);
   U276 : NAND2_X1 port map( A1 => n197, A2 => n39, ZN => n193);
   U277 : INV_X1 port map( A => n208, ZN => n197);
   U278 : XNOR2_X1 port map( A => n211, B => n210, ZN => SUM(15));
   U279 : OAI21_X1 port map( B1 => n22, B2 => n212, A => n189, ZN => n211);
   U280 : INV_X1 port map( A => n200, ZN => n212);
   U281 : INV_X1 port map( A => n5, ZN => n218);
   U282 : INV_X1 port map( A => n205, ZN => n196);
   U283 : XNOR2_X1 port map( A => n228, B => n229, ZN => SUM(11));
   U284 : OAI21_X1 port map( B1 => n230, B2 => n231, A => n226, ZN => n229);
   U285 : INV_X1 port map( A => n223, ZN => n231);
   U286 : INV_X1 port map( A => n232, ZN => n230);
   U287 : INV_X1 port map( A => n207, ZN => n238);
   U288 : INV_X1 port map( A => n163, ZN => n243);
   U289 : INV_X1 port map( A => n247, ZN => n246);
   U290 : INV_X1 port map( A => n253, ZN => n165);
   U291 : INV_X1 port map( A => n251, ZN => n254);
   U292 : INV_X1 port map( A => n44, ZN => n235);
   U293 : INV_X1 port map( A => n259, ZN => n258);
   U294 : INV_X1 port map( A => n261, ZN => n198);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_REGISTER_FILE_WINDOWING.all;

entity REGISTER_FILE_WINDOWING_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end REGISTER_FILE_WINDOWING_DW01_cmp6_0;

architecture SYN_rpl of REGISTER_FILE_WINDOWING_DW01_cmp6_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188 : std_logic;

begin
   
   U55 : NAND3_X1 port map( A1 => n76, A2 => n56, A3 => n57, ZN => n75);
   U57 : NAND3_X1 port map( A1 => n78, A2 => n54, A3 => n55, ZN => n77);
   U65 : NAND3_X1 port map( A1 => n89, A2 => n90, A3 => n91, ZN => n88);
   U67 : NAND3_X1 port map( A1 => n95, A2 => n93, A3 => n94, ZN => n92);
   U69 : NAND3_X1 port map( A1 => n97, A2 => n98, A3 => n99, ZN => n96);
   U73 : NAND3_X1 port map( A1 => n105, A2 => n64, A3 => n106, ZN => n104);
   U1 : OR2_X1 port map( A1 => A(12), A2 => n173, ZN => n150);
   U2 : AND2_X1 port map( A1 => B(31), A2 => n154, ZN => n63);
   U3 : AND2_X1 port map( A1 => n82, A2 => n51, ZN => n110);
   U4 : AND2_X1 port map( A1 => n85, A2 => n86, ZN => n111);
   U5 : AND2_X1 port map( A1 => n151, A2 => n150, ZN => n112);
   U6 : AND2_X1 port map( A1 => n149, A2 => n148, ZN => n113);
   U7 : AND2_X1 port map( A1 => n53, A2 => n52, ZN => n114);
   U8 : AND2_X1 port map( A1 => n139, A2 => n138, ZN => n115);
   U9 : AND2_X1 port map( A1 => n58, A2 => n48, ZN => n116);
   U10 : AND2_X1 port map( A1 => n137, A2 => n136, ZN => n117);
   U11 : AND2_X1 port map( A1 => n46, A2 => n47, ZN => n118);
   U12 : AND2_X1 port map( A1 => n147, A2 => n146, ZN => n119);
   U13 : CLKBUF_X1 port map( A => n175, Z => n120);
   U14 : OR2_X1 port map( A1 => B(1), A2 => n108, ZN => n121);
   U15 : OR2_X1 port map( A1 => n109, A2 => n186, ZN => n122);
   U16 : NAND3_X1 port map( A1 => n121, A2 => n122, A3 => n65, ZN => n107);
   U17 : OR2_X1 port map( A1 => A(8), A2 => n177, ZN => n123);
   U18 : OR2_X1 port map( A1 => A(9), A2 => n176, ZN => n124);
   U19 : NAND3_X1 port map( A1 => n96, A2 => n124, A3 => n123, ZN => n95);
   U20 : NAND2_X1 port map( A1 => n87, A2 => n111, ZN => n84);
   U21 : NAND2_X1 port map( A1 => n45, A2 => n43, ZN => n125);
   U22 : NAND2_X1 port map( A1 => n83, A2 => n110, ZN => n81);
   U23 : AND2_X1 port map( A1 => n141, A2 => n140, ZN => n126);
   U24 : AND2_X1 port map( A1 => n45, A2 => n43, ZN => n127);
   U25 : AND2_X1 port map( A1 => n118, A2 => n127, ZN => n131);
   U26 : NAND2_X1 port map( A1 => n129, A2 => n128, ZN => n68);
   U27 : AND2_X1 port map( A1 => n130, A2 => n126, ZN => n128);
   U28 : NAND2_X1 port map( A1 => n72, A2 => n131, ZN => n129);
   U29 : OR2_X1 port map( A1 => n125, A2 => n113, ZN => n130);
   U30 : AND2_X1 port map( A1 => n103, A2 => n102, ZN => n132);
   U31 : NAND2_X1 port map( A1 => n77, A2 => n115, ZN => n76);
   U32 : NAND2_X1 port map( A1 => n81, A2 => n117, ZN => n80);
   U33 : NOR2_X1 port map( A1 => n134, A2 => n135, ZN => n133);
   U34 : NOR2_X1 port map( A1 => n166, A2 => A(19), ZN => n134);
   U35 : NOR2_X1 port map( A1 => A(18), A2 => n167, ZN => n135);
   U36 : NAND2_X1 port map( A1 => n79, A2 => n133, ZN => n78);
   U37 : NAND2_X1 port map( A1 => n73, A2 => n119, ZN => n72);
   U38 : NAND2_X1 port map( A1 => n132, A2 => n101, ZN => n100);
   U39 : NAND2_X1 port map( A1 => n74, A2 => n116, ZN => n73);
   U40 : NAND2_X1 port map( A1 => n80, A2 => n114, ZN => n79);
   U41 : NAND2_X1 port map( A1 => n88, A2 => n112, ZN => n87);
   U42 : OR2_X1 port map( A1 => A(16), A2 => n169, ZN => n136);
   U43 : OR2_X1 port map( A1 => A(17), A2 => n168, ZN => n137);
   U44 : OR2_X1 port map( A1 => A(20), A2 => n165, ZN => n138);
   U45 : OR2_X1 port map( A1 => A(21), A2 => n164, ZN => n139);
   U46 : OR2_X1 port map( A1 => n157, A2 => A(28), ZN => n140);
   U47 : OR2_X1 port map( A1 => A(29), A2 => n156, ZN => n141);
   U48 : OR2_X1 port map( A1 => A(14), A2 => n171, ZN => n142);
   U49 : OR2_X1 port map( A1 => n170, A2 => A(15), ZN => n143);
   U50 : NAND3_X1 port map( A1 => n84, A2 => n143, A3 => n142, ZN => n83);
   U51 : OR2_X1 port map( A1 => A(22), A2 => n163, ZN => n144);
   U52 : OR2_X1 port map( A1 => A(23), A2 => n162, ZN => n145);
   U53 : NAND3_X1 port map( A1 => n144, A2 => n145, A3 => n75, ZN => n74);
   U54 : OR2_X1 port map( A1 => A(24), A2 => n161, ZN => n146);
   U56 : OR2_X1 port map( A1 => A(25), A2 => n160, ZN => n147);
   U58 : OR2_X1 port map( A1 => A(26), A2 => n159, ZN => n148);
   U59 : OR2_X1 port map( A1 => n158, A2 => A(27), ZN => n149);
   U60 : OR2_X1 port map( A1 => n172, A2 => A(13), ZN => n151);
   U61 : OAI22_X1 port map( A1 => B(31), A2 => n154, B1 => n63, B2 => n66, ZN 
                           => n152);
   U62 : INV_X1 port map( A => A(30), ZN => n155);
   U63 : NAND2_X1 port map( A1 => A(18), A2 => n167, ZN => n53);
   U64 : NAND2_X1 port map( A1 => A(19), A2 => n166, ZN => n54);
   U66 : NAND2_X1 port map( A1 => A(9), A2 => n176, ZN => n94);
   U68 : OR2_X1 port map( A1 => n155, A2 => B(30), ZN => n42);
   U70 : NAND2_X1 port map( A1 => A(5), A2 => n180, ZN => n102);
   U71 : NOR4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => EQ
                           );
   U72 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n37);
   U74 : NAND2_X1 port map( A1 => A(12), A2 => n173, ZN => n89);
   U75 : NAND2_X1 port map( A1 => A(17), A2 => n168, ZN => n52);
   U76 : NAND2_X1 port map( A1 => A(29), A2 => n156, ZN => n41);
   U77 : NAND2_X1 port map( A1 => A(20), A2 => n165, ZN => n55);
   U78 : INV_X1 port map( A => A(1), ZN => n186);
   U79 : NAND4_X1 port map( A1 => n45, A2 => n46, A3 => n47, A4 => n48, ZN => 
                           n38);
   U80 : AND4_X1 port map( A1 => n51, A2 => n52, A3 => n53, A4 => n54, ZN => 
                           n50);
   U81 : INV_X1 port map( A => A(31), ZN => n154);
   U82 : AND2_X1 port map( A1 => n42, A2 => n41, ZN => n67);
   U83 : OAI221_X1 port map( B1 => A(4), B2 => n181, C1 => A(5), C2 => n180, A 
                           => n104, ZN => n103);
   U84 : NAND2_X1 port map( A1 => A(4), A2 => n181, ZN => n105);
   U85 : AND2_X1 port map( A1 => n186, A2 => n109, ZN => n108);
   U86 : NOR2_X1 port map( A1 => n188, A2 => A(0), ZN => n109);
   U87 : NAND2_X1 port map( A1 => A(2), A2 => n185, ZN => n65);
   U88 : INV_X1 port map( A => B(18), ZN => n167);
   U89 : NAND2_X1 port map( A1 => A(8), A2 => n177, ZN => n97);
   U90 : NAND2_X1 port map( A1 => A(13), A2 => n172, ZN => n86);
   U91 : INV_X1 port map( A => B(19), ZN => n166);
   U92 : INV_X1 port map( A => B(5), ZN => n180);
   U93 : INV_X1 port map( A => B(9), ZN => n176);
   U94 : NAND2_X1 port map( A1 => A(22), A2 => n163, ZN => n57);
   U95 : NAND2_X1 port map( A1 => A(3), A2 => n183, ZN => n64);
   U96 : NOR4_X1 port map( A1 => n152, A2 => n63, A3 => n184, A4 => n182, ZN =>
                           n62);
   U97 : INV_X1 port map( A => n65, ZN => n184);
   U98 : INV_X1 port map( A => n64, ZN => n182);
   U99 : NAND2_X1 port map( A1 => A(26), A2 => n159, ZN => n46);
   U100 : INV_X1 port map( A => B(12), ZN => n173);
   U101 : NAND2_X1 port map( A1 => A(23), A2 => n162, ZN => n58);
   U102 : NAND2_X1 port map( A1 => A(27), A2 => n158, ZN => n45);
   U103 : INV_X1 port map( A => B(17), ZN => n168);
   U104 : INV_X1 port map( A => B(29), ZN => n156);
   U105 : NAND2_X1 port map( A1 => A(28), A2 => n157, ZN => n43);
   U106 : NAND2_X1 port map( A1 => A(16), A2 => n169, ZN => n51);
   U107 : NAND2_X1 port map( A1 => A(25), A2 => n160, ZN => n47);
   U108 : INV_X1 port map( A => B(20), ZN => n165);
   U109 : NAND2_X1 port map( A1 => A(21), A2 => n164, ZN => n56);
   U110 : NAND2_X1 port map( A1 => A(24), A2 => n161, ZN => n48);
   U111 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n39);
   U112 : OAI22_X1 port map( A1 => A(1), A2 => n44, B1 => n44, B2 => n187, ZN 
                           => n40);
   U113 : AND2_X1 port map( A1 => A(0), A2 => n188, ZN => n44);
   U114 : INV_X1 port map( A => B(1), ZN => n187);
   U115 : INV_X1 port map( A => B(8), ZN => n177);
   U116 : INV_X1 port map( A => B(13), ZN => n172);
   U117 : INV_X1 port map( A => B(22), ZN => n163);
   U118 : INV_X1 port map( A => B(3), ZN => n183);
   U119 : INV_X1 port map( A => B(26), ZN => n159);
   U120 : INV_X1 port map( A => B(23), ZN => n162);
   U121 : INV_X1 port map( A => B(27), ZN => n158);
   U122 : INV_X1 port map( A => B(0), ZN => n188);
   U123 : INV_X1 port map( A => B(28), ZN => n157);
   U124 : INV_X1 port map( A => B(16), ZN => n169);
   U125 : INV_X1 port map( A => B(25), ZN => n160);
   U126 : INV_X1 port map( A => B(21), ZN => n164);
   U127 : INV_X1 port map( A => B(24), ZN => n161);
   U128 : INV_X1 port map( A => B(4), ZN => n181);
   U129 : OAI22_X1 port map( A1 => B(31), A2 => n154, B1 => n66, B2 => n63, ZN 
                           => LT);
   U130 : AND4_X1 port map( A1 => n55, A2 => n56, A3 => n57, A4 => n58, ZN => 
                           n49);
   U131 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           n36);
   U132 : INV_X1 port map( A => B(2), ZN => n185);
   U133 : OAI221_X1 port map( B1 => A(2), B2 => n185, C1 => A(3), C2 => n183, A
                           => n107, ZN => n106);
   U134 : NAND2_X1 port map( A1 => A(7), A2 => n178, ZN => n98);
   U135 : NAND2_X1 port map( A1 => A(11), A2 => n174, ZN => n90);
   U136 : INV_X1 port map( A => B(11), ZN => n174);
   U137 : AND4_X1 port map( A1 => n105, A2 => n102, A3 => n101, A4 => n98, ZN 
                           => n61);
   U138 : INV_X1 port map( A => B(7), ZN => n178);
   U139 : AND4_X1 port map( A1 => n89, A2 => n86, A3 => n85, A4 => n82, ZN => 
                           n59);
   U140 : NAND2_X1 port map( A1 => n170, A2 => A(15), ZN => n82);
   U141 : AND4_X1 port map( A1 => n97, A2 => n94, A3 => n93, A4 => n90, ZN => 
                           n60);
   U142 : OAI221_X1 port map( B1 => A(10), B2 => n120, C1 => n174, C2 => A(11),
                           A => n92, ZN => n91);
   U143 : NAND2_X1 port map( A1 => n175, A2 => A(10), ZN => n93);
   U144 : OAI221_X1 port map( B1 => A(6), B2 => n179, C1 => n178, C2 => A(7), A
                           => n100, ZN => n99);
   U145 : NAND2_X1 port map( A1 => A(6), A2 => n179, ZN => n101);
   U146 : NAND2_X1 port map( A1 => n171, A2 => A(14), ZN => n85);
   U147 : INV_X1 port map( A => B(10), ZN => n175);
   U148 : INV_X1 port map( A => B(6), ZN => n179);
   U149 : INV_X1 port map( A => B(14), ZN => n171);
   U150 : INV_X1 port map( A => B(15), ZN => n170);
   U151 : AOI22_X1 port map( A1 => B(30), A2 => n155, B1 => n68, B2 => n67, ZN 
                           => n66);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_REGISTER_FILE_WINDOWING.all;

entity REGISTER_FILE_WINDOWING_DW01_addsub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in std_logic;
         SUM : out std_logic_vector (31 downto 0);  CO : out std_logic);

end REGISTER_FILE_WINDOWING_DW01_addsub_0;

architecture SYN_rpl of REGISTER_FILE_WINDOWING_DW01_addsub_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n63 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => A(30), B => n32, Z => SUM(30));
   U3 : XOR2_X1 port map( A => A(29), B => n33, Z => SUM(29));
   U4 : XOR2_X1 port map( A => A(28), B => n34, Z => SUM(28));
   U5 : XOR2_X1 port map( A => A(27), B => n35, Z => SUM(27));
   U6 : XOR2_X1 port map( A => A(26), B => n36, Z => SUM(26));
   U7 : XOR2_X1 port map( A => A(25), B => n37, Z => SUM(25));
   U8 : XOR2_X1 port map( A => A(24), B => n38, Z => SUM(24));
   U9 : XOR2_X1 port map( A => A(23), B => n39, Z => SUM(23));
   U10 : XOR2_X1 port map( A => A(22), B => n40, Z => SUM(22));
   U11 : XOR2_X1 port map( A => A(21), B => n41, Z => SUM(21));
   U12 : XOR2_X1 port map( A => A(20), B => n42, Z => SUM(20));
   U13 : XOR2_X1 port map( A => A(19), B => n43, Z => SUM(19));
   U14 : XOR2_X1 port map( A => A(18), B => n44, Z => SUM(18));
   U15 : XOR2_X1 port map( A => A(17), B => n45, Z => SUM(17));
   U16 : XOR2_X1 port map( A => A(16), B => n46, Z => SUM(16));
   U17 : XOR2_X1 port map( A => A(15), B => n47, Z => SUM(15));
   U18 : XOR2_X1 port map( A => A(14), B => n48, Z => SUM(14));
   U19 : XOR2_X1 port map( A => A(13), B => n49, Z => SUM(13));
   U20 : XOR2_X1 port map( A => A(12), B => n50, Z => SUM(12));
   U21 : XOR2_X1 port map( A => A(11), B => n51, Z => SUM(11));
   U22 : XOR2_X1 port map( A => A(10), B => n52, Z => SUM(10));
   U23 : XOR2_X1 port map( A => A(9), B => n53, Z => SUM(9));
   U24 : XOR2_X1 port map( A => A(8), B => n54, Z => SUM(8));
   U25 : XOR2_X1 port map( A => A(7), B => n55, Z => SUM(7));
   U26 : XOR2_X1 port map( A => A(6), B => n56, Z => SUM(6));
   U27 : XOR2_X1 port map( A => A(5), B => n57, Z => SUM(5));
   U28 : XOR2_X1 port map( A => A(4), B => n58, Z => SUM(4));
   U29 : XOR2_X1 port map( A => A(3), B => n59, Z => SUM(3));
   U30 : XOR2_X1 port map( A => A(2), B => n60, Z => SUM(2));
   U32 : XOR2_X1 port map( A => A(1), B => A(0), Z => SUM(1));
   U1 : XNOR2_X1 port map( A => A(31), B => n63, ZN => SUM(31));
   U31 : NAND2_X1 port map( A1 => A(30), A2 => n32, ZN => n63);
   U33 : AND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n60);
   U34 : AND2_X1 port map( A1 => A(4), A2 => n58, ZN => n57);
   U35 : AND2_X1 port map( A1 => A(8), A2 => n54, ZN => n53);
   U36 : AND2_X1 port map( A1 => A(9), A2 => n53, ZN => n52);
   U37 : AND2_X1 port map( A1 => A(19), A2 => n43, ZN => n42);
   U38 : AND2_X1 port map( A1 => A(20), A2 => n42, ZN => n41);
   U39 : AND2_X1 port map( A1 => A(21), A2 => n41, ZN => n40);
   U40 : AND2_X1 port map( A1 => A(2), A2 => n60, ZN => n59);
   U41 : AND2_X1 port map( A1 => A(3), A2 => n59, ZN => n58);
   U42 : AND2_X1 port map( A1 => A(5), A2 => n57, ZN => n56);
   U43 : AND2_X1 port map( A1 => A(6), A2 => n56, ZN => n55);
   U44 : AND2_X1 port map( A1 => A(7), A2 => n55, ZN => n54);
   U45 : AND2_X1 port map( A1 => A(10), A2 => n52, ZN => n51);
   U46 : AND2_X1 port map( A1 => A(11), A2 => n51, ZN => n50);
   U47 : AND2_X1 port map( A1 => A(12), A2 => n50, ZN => n49);
   U48 : AND2_X1 port map( A1 => A(13), A2 => n49, ZN => n48);
   U49 : AND2_X1 port map( A1 => A(14), A2 => n48, ZN => n47);
   U50 : AND2_X1 port map( A1 => A(15), A2 => n47, ZN => n46);
   U51 : AND2_X1 port map( A1 => A(16), A2 => n46, ZN => n45);
   U52 : AND2_X1 port map( A1 => A(17), A2 => n45, ZN => n44);
   U53 : AND2_X1 port map( A1 => A(18), A2 => n44, ZN => n43);
   U54 : AND2_X1 port map( A1 => A(22), A2 => n40, ZN => n39);
   U55 : AND2_X1 port map( A1 => A(23), A2 => n39, ZN => n38);
   U56 : AND2_X1 port map( A1 => A(24), A2 => n38, ZN => n37);
   U57 : AND2_X1 port map( A1 => A(25), A2 => n37, ZN => n36);
   U58 : AND2_X1 port map( A1 => A(26), A2 => n36, ZN => n35);
   U59 : AND2_X1 port map( A1 => A(27), A2 => n35, ZN => n34);
   U60 : AND2_X1 port map( A1 => A(28), A2 => n34, ZN => n33);
   U61 : AND2_X1 port map( A1 => A(29), A2 => n33, ZN => n32);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_REGISTER_FILE_WINDOWING.all;

entity REGISTER_FILE_WINDOWING is

   port( CLK, RESET, ENABLE, RD1, RD2, WR, CALL, SIGRETURN : in std_logic;  
         ADD_WR, ADD_RD1, ADD_RD2 : in std_logic_vector (3 downto 0);  DATAIN :
         in std_logic_vector (63 downto 0);  OUT1, OUT2, MEM_BUS : out 
         std_logic_vector (63 downto 0);  MEM_BUSread : in std_logic_vector (63
         downto 0);  FILL, SPILL : out std_logic);

end REGISTER_FILE_WINDOWING;

architecture SYN_BEHAVIORAL of REGISTER_FILE_WINDOWING is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component REGISTER_FILE_WINDOWING_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component REGISTER_FILE_WINDOWING_DW01_addsub_2
      port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (31 downto 0);  CO : out 
            std_logic);
   end component;
   
   component REGISTER_FILE_WINDOWING_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component REGISTER_FILE_WINDOWING_DW01_addsub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI, ADD_SUB : in 
            std_logic;  SUM : out std_logic_vector (31 downto 0);  CO : out 
            std_logic);
   end component;
   
   signal OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, OUT1_59_port,
      OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, OUT1_54_port, 
      OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, OUT1_49_port, 
      OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, OUT1_44_port, 
      OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, OUT1_39_port, 
      OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, OUT1_34_port, 
      OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, OUT1_29_port, 
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, MEM_BUS_63_port, 
      MEM_BUS_62_port, MEM_BUS_61_port, MEM_BUS_60_port, MEM_BUS_59_port, 
      MEM_BUS_58_port, MEM_BUS_57_port, MEM_BUS_56_port, MEM_BUS_55_port, 
      MEM_BUS_54_port, MEM_BUS_53_port, MEM_BUS_52_port, MEM_BUS_51_port, 
      MEM_BUS_50_port, MEM_BUS_49_port, MEM_BUS_48_port, MEM_BUS_47_port, 
      MEM_BUS_46_port, MEM_BUS_45_port, MEM_BUS_44_port, MEM_BUS_43_port, 
      MEM_BUS_42_port, MEM_BUS_41_port, MEM_BUS_40_port, MEM_BUS_39_port, 
      MEM_BUS_38_port, MEM_BUS_37_port, MEM_BUS_36_port, MEM_BUS_35_port, 
      MEM_BUS_34_port, MEM_BUS_33_port, MEM_BUS_32_port, MEM_BUS_31_port, 
      MEM_BUS_30_port, MEM_BUS_29_port, MEM_BUS_28_port, MEM_BUS_27_port, 
      MEM_BUS_26_port, MEM_BUS_25_port, MEM_BUS_24_port, MEM_BUS_23_port, 
      MEM_BUS_22_port, MEM_BUS_21_port, MEM_BUS_20_port, MEM_BUS_19_port, 
      MEM_BUS_18_port, MEM_BUS_17_port, MEM_BUS_16_port, MEM_BUS_15_port, 
      MEM_BUS_14_port, MEM_BUS_13_port, MEM_BUS_12_port, MEM_BUS_11_port, 
      MEM_BUS_10_port, MEM_BUS_9_port, MEM_BUS_8_port, MEM_BUS_7_port, 
      MEM_BUS_6_port, MEM_BUS_5_port, MEM_BUS_4_port, MEM_BUS_3_port, 
      MEM_BUS_2_port, MEM_BUS_1_port, MEM_BUS_0_port, CWP_31_port, CWP_30_port,
      CWP_29_port, CWP_28_port, CWP_27_port, CWP_26_port, CWP_25_port, 
      CWP_24_port, CWP_23_port, CWP_22_port, CWP_21_port, CWP_20_port, 
      CWP_19_port, CWP_18_port, CWP_17_port, CWP_16_port, CWP_15_port, 
      CWP_14_port, CWP_13_port, CWP_12_port, CWP_11_port, CWP_10_port, 
      CWP_9_port, CWP_8_port, CWP_7_port, CWP_6_port, CWP_5_port, CWP_4_port, 
      CWP_3_port, CWP_2_port, CWP_1_port, CWP_0_port, N75, N76, N77, N78, N79, 
      N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94
      , N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N139
      , N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
      N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
      N234, N235, N236, N237, N238, N239, N240, N241, i_31_port, i_30_port, 
      i_29_port, i_28_port, i_27_port, i_26_port, i_25_port, i_24_port, 
      i_23_port, i_22_port, i_21_port, i_20_port, i_19_port, i_18_port, 
      i_17_port, i_16_port, i_15_port, i_14_port, i_13_port, i_12_port, 
      i_11_port, i_10_port, i_9_port, i_8_port, i_7_port, i_6_port, i_5_port, 
      i_4_port, i_3_port, i_2_port, i_1_port, i_0_port, N623, N624, N625, N626,
      N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, 
      N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, 
      N651, N652, N653, N2739, U3_U1_Z_0, U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3, 
      U3_U1_Z_4, U3_U1_Z_5, U3_U1_Z_6, U3_U1_Z_7, U3_U1_Z_8, U3_U1_Z_9, 
      U3_U1_Z_10, U3_U1_Z_11, U3_U1_Z_12, U3_U1_Z_13, U3_U1_Z_14, U3_U1_Z_15, 
      U3_U1_Z_16, U3_U1_Z_17, U3_U1_Z_18, U3_U1_Z_19, U3_U1_Z_20, U3_U1_Z_21, 
      U3_U1_Z_22, U3_U1_Z_23, U3_U1_Z_24, U3_U1_Z_25, U3_U1_Z_26, U3_U1_Z_27, 
      U3_U1_Z_28, U3_U1_Z_29, U3_U1_Z_30, U3_U1_Z_31, U3_U2_Z_0, U3_U2_Z_1, 
      U3_U2_Z_2, U3_U2_Z_3, U3_U2_Z_4, U3_U2_Z_5, U3_U2_Z_6, U3_U2_Z_7, 
      U3_U2_Z_8, U3_U2_Z_9, U3_U2_Z_10, U3_U2_Z_11, U3_U2_Z_12, U3_U2_Z_13, 
      U3_U2_Z_14, U3_U2_Z_15, U3_U2_Z_16, U3_U2_Z_17, U3_U2_Z_18, U3_U2_Z_19, 
      U3_U2_Z_20, U3_U2_Z_21, U3_U2_Z_22, U3_U2_Z_23, U3_U2_Z_24, U3_U2_Z_25, 
      U3_U2_Z_26, U3_U2_Z_27, U3_U2_Z_28, U3_U2_Z_29, U3_U2_Z_30, U3_U2_Z_31, 
      U3_U3_Z_0, U3_U3_Z_1, U3_U3_Z_2, U3_U3_Z_3, U3_U3_Z_4, U3_U3_Z_5, 
      U3_U3_Z_6, U3_U3_Z_7, U3_U3_Z_8, U3_U3_Z_9, U3_U3_Z_10, U3_U3_Z_11, 
      U3_U3_Z_12, U3_U3_Z_13, U3_U3_Z_14, U3_U3_Z_15, U3_U3_Z_16, U3_U3_Z_17, 
      U3_U3_Z_18, U3_U3_Z_19, U3_U3_Z_20, U3_U3_Z_21, U3_U3_Z_22, U3_U3_Z_23, 
      U3_U3_Z_24, U3_U3_Z_25, U3_U3_Z_26, U3_U3_Z_27, U3_U3_Z_28, U3_U3_Z_29, 
      U3_U3_Z_30, U3_U3_Z_31, U3_U7_Z_0, U3_U7_Z_1, U3_U7_Z_2, U3_U7_Z_3, 
      U3_U7_Z_4, U3_U7_Z_5, U3_U7_Z_6, U3_U7_Z_7, U3_U7_Z_8, U3_U7_Z_9, 
      U3_U7_Z_10, U3_U7_Z_11, U3_U7_Z_12, U3_U7_Z_13, U3_U7_Z_14, U3_U7_Z_15, 
      U3_U7_Z_16, U3_U7_Z_17, U3_U7_Z_18, U3_U7_Z_19, U3_U7_Z_20, U3_U7_Z_21, 
      U3_U7_Z_22, U3_U7_Z_23, U3_U7_Z_24, U3_U7_Z_25, U3_U7_Z_26, U3_U7_Z_27, 
      U3_U7_Z_28, U3_U7_Z_29, U3_U7_Z_30, U3_U7_Z_31, U3_U8_Z_0, U3_U8_Z_2, 
      U3_U8_Z_3, U3_U9_Z_0, n967, n968, n969, n970, n971, n972, n973, n974, 
      n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, 
      n987, n988, n989, n990, n991, n992, n993, n994, n3043, n3044, n3045, 
      n3046, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, 
      n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, 
      n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, 
      n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, 
      n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
      n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, 
      n3136, n3137, n3138, n3139, n3140, n3141, n3236, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, 
      n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, 
      n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, 
      n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, 
      n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, 
      n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, 
      n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, 
      n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, 
      n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, 
      n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, 
      n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, 
      n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, 
      n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, 
      n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, 
      n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, 
      n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, 
      n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, 
      n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, 
      n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, 
      n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, 
      n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, 
      n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, 
      n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, 
      n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, 
      n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, 
      n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, 
      n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, 
      n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, 
      n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, 
      n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
      n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, 
      n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, 
      n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, 
      n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, 
      n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, 
      n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
      n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, 
      n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
      n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, 
      n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
      n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, 
      n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
      n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, 
      n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
      n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
      n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, 
      n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
      n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
      n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, 
      n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
      n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
      n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
      n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, 
      n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
      n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, 
      n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
      n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, 
      n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
      n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, 
      n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
      n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, 
      n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, 
      n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
      n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, 
      n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, 
      n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, 
      n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, 
      n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, 
      n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, 
      n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, 
      n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, 
      n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, 
      n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, 
      n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, 
      n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, 
      n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, 
      n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, 
      n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, 
      n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, 
      n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, 
      n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, 
      n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, 
      n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, 
      n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, 
      n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, 
      n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, 
      n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, 
      n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, 
      n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
      n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
      n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
      n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, 
      n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, 
      n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, 
      n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, 
      n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, 
      n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
      n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, 
      n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, 
      n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
      n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, 
      n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, 
      n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, 
      n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, 
      n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, 
      n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, 
      n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, 
      n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, 
      n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, 
      n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, 
      n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, 
      n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, 
      n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, 
      n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, 
      n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, 
      n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, 
      n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, 
      n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, 
      n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, 
      n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, 
      n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, 
      n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, 
      n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, 
      n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, 
      n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, 
      n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, 
      n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, 
      n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, 
      n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, 
      n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, 
      n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, 
      n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, 
      n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, 
      n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, 
      n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, 
      n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, 
      n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, 
      n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, 
      n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, 
      n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, 
      n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, 
      n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, 
      n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, 
      n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, 
      n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, 
      n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, 
      n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, 
      n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, 
      n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, 
      n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, 
      n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, 
      n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, 
      n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, 
      n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, 
      n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, 
      n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, 
      n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, 
      n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, 
      n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, 
      n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, 
      n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, 
      n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, 
      n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, 
      n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, 
      n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, 
      n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, 
      n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, 
      n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, 
      n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, 
      n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, 
      n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, 
      n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, 
      n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, 
      n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, 
      n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, 
      n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, 
      n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, 
      n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, 
      n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, 
      n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5609, n5610, n5611, 
      n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
      n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
      n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5699, n5700, n5731, n5732, n5733, n5734, 
      n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, 
      n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, 
      n5755, n5756, n13211, n13212, n13213, n13214, n13215, n13216, n13217, 
      n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, 
      n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, 
      n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, 
      n13245, n13246, n13247, n13248, n15107, n15108, n15109, n15110, n15111, 
      n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, 
      n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, 
      n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, 
      n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, 
      n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, 
      n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, 
      n15166, n15167, n15168, n15169, n15170, n15175, n15176, n15178, n15179, 
      n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, 
      n15189, n15190, n15191, n15192, n15193, n15194, n15197, n15200, n15201, 
      n15202, n15203, n15204, n15205, n15207, n15208, n15210, n15211, n15212, 
      n15213, n15214, n15215, n15216, n15217, n15218, n15220, n15221, n15222, 
      n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, 
      n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, 
      n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, 
      n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, 
      n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, 
      n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, 
      n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, 
      n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, 
      n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, 
      n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, 
      n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, 
      n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, 
      n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, 
      n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, 
      n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, 
      n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, 
      n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, 
      n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, 
      n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, 
      n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, 
      n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, 
      n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, 
      n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, 
      n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, 
      n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, 
      n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, 
      n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, 
      n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, 
      n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, 
      n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, 
      n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, 
      n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, 
      n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, 
      n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, 
      n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, 
      n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, 
      n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, 
      n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, 
      n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, 
      n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, 
      n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, 
      n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, 
      n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, 
      n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, 
      n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, 
      n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, 
      n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, 
      n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, 
      n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, 
      n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, 
      n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, 
      n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, 
      n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, 
      n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, 
      n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, 
      n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, 
      n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, 
      n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, 
      n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, 
      n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, 
      n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, 
      n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, 
      n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, 
      n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, 
      n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, 
      n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, 
      n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, 
      n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, 
      n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, 
      n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, 
      n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, 
      n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, 
      n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, 
      n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, 
      n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, 
      n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, 
      n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, 
      n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, 
      n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, 
      n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, 
      n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, 
      n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, 
      n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, 
      n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, 
      n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, 
      n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, 
      n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, 
      n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, 
      n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, 
      n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, 
      n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, 
      n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, 
      n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, 
      n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, 
      n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, 
      n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, 
      n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, 
      n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, 
      n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, 
      n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, 
      n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, 
      n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, 
      n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, 
      n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, 
      n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, 
      n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, 
      n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, 
      n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, 
      n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, 
      n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, 
      n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, 
      n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, 
      n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, 
      n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, 
      n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, 
      n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, 
      n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, 
      n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, 
      n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, 
      n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, 
      n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, 
      n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, 
      n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, 
      n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, 
      n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, 
      n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, 
      n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, 
      n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, 
      n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, 
      n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, 
      n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, 
      n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, 
      n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, 
      n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, 
      n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, 
      n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, 
      n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, 
      n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, 
      n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, 
      n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, 
      n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, 
      n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, 
      n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, 
      n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, 
      n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, 
      n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, 
      n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, 
      n16546, n16549, n16552, n16553, n16554, n16555, n16579, n16580, n16581, 
      n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, 
      n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, 
      n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, 
      n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, 
      n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, 
      n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, 
      n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, 
      n16664, n16668, n16673, n16678, n16683, n16713, n16716, n16718, n16719, 
      n16720, n16721, n16722, n16724, n16725, n16728, n16730, n16731, n16732, 
      n16733, n16734, n16735, n16770, n16771, n16774, n16775, n16779, n16784, 
      n16787, n16788, n16790, n16791, n16795, n16796, n16802, n16823, n16824, 
      n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, 
      n16836, n16850, n16851, n16854, n16855, n16856, n16857, n16858, n16859, 
      n16860, n16861, n16862, n16863, n16877, n16878, n16881, n16882, n16883, 
      n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16904, n16905, 
      n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, 
      n16917, n16931, n16932, n16935, n16936, n16937, n16938, n16939, n16940, 
      n16941, n16942, n16943, n16944, n16958, n16959, n16962, n16963, n16964, 
      n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16985, n16986, 
      n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, 
      n16998, n17012, n17013, n17016, n17017, n17018, n17019, n17020, n17021, 
      n17022, n17023, n17024, n17025, n17039, n17040, n17043, n17044, n17045, 
      n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17066, n17067, 
      n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, 
      n17079, n17093, n17094, n17097, n17098, n17099, n17100, n17101, n17102, 
      n17103, n17104, n17105, n17106, n17120, n17121, n17124, n17125, n17126, 
      n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17147, n17148, 
      n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, 
      n17160, n17174, n17175, n17178, n17179, n17180, n17181, n17182, n17183, 
      n17184, n17185, n17186, n17187, n17201, n17202, n17205, n17206, n17207, 
      n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17228, n17229, 
      n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, 
      n17241, n17255, n17256, n17259, n17260, n17261, n17262, n17263, n17264, 
      n17265, n17266, n17267, n17268, n17282, n17283, n17286, n17287, n17288, 
      n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17309, n17310, 
      n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, 
      n17322, n17336, n17337, n17340, n17341, n17342, n17343, n17344, n17345, 
      n17346, n17347, n17348, n17349, n17363, n17364, n17367, n17368, n17369, 
      n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17390, n17391, 
      n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, 
      n17403, n17417, n17418, n17421, n17422, n17423, n17424, n17425, n17426, 
      n17427, n17428, n17429, n17430, n17444, n17445, n17448, n17449, n17450, 
      n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17471, n17472, 
      n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, 
      n17484, n17498, n17499, n17502, n17503, n17504, n17505, n17506, n17507, 
      n17508, n17509, n17510, n17511, n17525, n17526, n17529, n17530, n17531, 
      n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17552, n17553, 
      n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, 
      n17565, n17579, n17580, n17583, n17584, n17585, n17586, n17587, n17588, 
      n17589, n17590, n17591, n17592, n17606, n17607, n17610, n17611, n17612, 
      n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17633, n17634, 
      n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, 
      n17646, n17660, n17661, n17664, n17665, n17666, n17667, n17668, n17669, 
      n17670, n17671, n17672, n17673, n17687, n17688, n17691, n17692, n17693, 
      n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17714, n17715, 
      n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, 
      n17727, n17741, n17742, n17745, n17746, n17747, n17748, n17749, n17750, 
      n17751, n17752, n17753, n17754, n17768, n17769, n17772, n17773, n17774, 
      n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17795, n17796, 
      n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, 
      n17808, n17822, n17823, n17826, n17827, n17828, n17829, n17830, n17831, 
      n17832, n17833, n17834, n17835, n17849, n17850, n17853, n17854, n17855, 
      n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17876, n17877, 
      n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, 
      n17889, n17903, n17904, n17907, n17908, n17909, n17910, n17911, n17912, 
      n17913, n17914, n17915, n17916, n17930, n17931, n17934, n17935, n17936, 
      n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17957, n17958, 
      n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, 
      n17970, n17984, n17985, n17988, n17989, n17990, n17991, n17992, n17993, 
      n17994, n17995, n17996, n17997, n18011, n18012, n18015, n18016, n18017, 
      n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18038, n18039, 
      n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, 
      n18051, n18065, n18066, n18069, n18070, n18071, n18072, n18073, n18074, 
      n18075, n18076, n18077, n18078, n18092, n18093, n18096, n18097, n18098, 
      n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18119, n18120, 
      n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, 
      n18132, n18146, n18147, n18150, n18151, n18152, n18153, n18154, n18155, 
      n18156, n18157, n18158, n18159, n18173, n18174, n18177, n18178, n18179, 
      n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18200, n18201, 
      n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, 
      n18213, n18227, n18228, n18231, n18232, n18233, n18234, n18235, n18236, 
      n18237, n18238, n18239, n18240, n18254, n18255, n18258, n18259, n18260, 
      n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18281, n18282, 
      n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, 
      n18294, n18308, n18309, n18312, n18313, n18314, n18315, n18316, n18317, 
      n18318, n18319, n18320, n18321, n18335, n18336, n18339, n18340, n18341, 
      n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18362, n18363, 
      n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, 
      n18375, n18389, n18390, n18393, n18394, n18395, n18396, n18397, n18398, 
      n18399, n18400, n18401, n18402, n18416, n18417, n18420, n18421, n18422, 
      n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18443, n18444, 
      n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, 
      n18456, n18470, n18471, n18474, n18475, n18476, n18477, n18478, n18479, 
      n18480, n18481, n18482, n18483, n18509, n18510, n18513, n18514, n18515, 
      n18516, n18517, n18518, n18519, n18520, n18522, n18523, n18525, n18526, 
      n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, 
      n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, 
      n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, 
      n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, 
      n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, 
      n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, 
      n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, 
      n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, 
      n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, 
      n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, 
      n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, 
      n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, 
      n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, 
      n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, 
      n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, 
      n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, 
      n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, 
      n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, 
      n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, 
      n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, 
      n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, 
      n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, 
      n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, 
      n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, 
      n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, 
      n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, 
      n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, 
      n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, 
      n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, 
      n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, 
      n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, 
      n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, 
      n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, 
      n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, 
      n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, 
      n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, 
      n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, 
      n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, 
      n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, 
      n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, 
      n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, 
      n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, 
      n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, 
      n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, 
      n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, 
      n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, 
      n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, 
      n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, 
      n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, 
      n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, 
      n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, 
      n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, 
      n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, 
      n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, 
      n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, 
      n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, 
      n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, 
      n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, 
      n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, 
      n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, 
      n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, 
      n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, 
      n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, 
      n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, 
      n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, 
      n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, 
      n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, 
      n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, 
      n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, 
      n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, 
      n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, 
      n19323, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, 
      n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, 
      n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, 
      n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, 
      n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, 
      n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, 
      n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, 
      n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, 
      n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, 
      n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, 
      n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, 
      n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, 
      n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, 
      n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, 
      n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, 
      n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, 
      n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, 
      n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, 
      n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, 
      n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, 
      n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, 
      n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, 
      n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, 
      n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, 
      n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, 
      n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, 
      n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, 
      n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, 
      n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, 
      n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, 
      n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, 
      n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, 
      n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, 
      n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, 
      n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, 
      n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, 
      n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, 
      n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, 
      n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, 
      n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, 
      n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, 
      n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, 
      n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, 
      n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, 
      n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, 
      n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, 
      n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, 
      n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, 
      n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, 
      n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, 
      n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, 
      n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, 
      n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, 
      n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, 
      n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, 
      n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, 
      n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, 
      n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, 
      n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, 
      n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, 
      n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, 
      n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, 
      n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, 
      n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, 
      n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, 
      n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, 
      n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, 
      n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, 
      n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, 
      n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, 
      n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, 
      n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, 
      n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, 
      n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, 
      n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, 
      n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, 
      n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, 
      n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, 
      n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, 
      n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, 
      n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, 
      n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, 
      n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, 
      n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, 
      n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, 
      n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, 
      n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, 
      n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, 
      n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, 
      n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, 
      n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, 
      n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, 
      n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, 
      n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, 
      n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, 
      n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, 
      n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, 
      n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, 
      n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, 
      n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, 
      n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, 
      n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, 
      n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, 
      n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, 
      n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, 
      n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, 
      n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, 
      n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, 
      n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, 
      n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, 
      n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, 
      n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, 
      n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, 
      n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, 
      n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, 
      n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, 
      n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, 
      n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, 
      n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, 
      n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, 
      n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, 
      n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, 
      n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, 
      n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, 
      n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, 
      n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, 
      n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, 
      n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, 
      n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, 
      n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, 
      n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, 
      n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, 
      n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, 
      n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, 
      n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, 
      n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, 
      n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, 
      n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, 
      n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, 
      n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, 
      n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, 
      n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, 
      n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, 
      n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, 
      n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, 
      n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, 
      n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, 
      n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, 
      n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, 
      n20728, n20729, n20730, n20731, n20732, n20734, n20736, n20750, n20752, 
      n20753, n20754, n20756, n20759, n20760, n20761, n20764, n20765, n20766, 
      n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, 
      n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, 
      n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, 
      n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, 
      n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, 
      n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, 
      n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, 
      n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, 
      n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, 
      n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, 
      n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, 
      n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, 
      n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, 
      n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, 
      n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, 
      n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, 
      n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, 
      n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, 
      n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, 
      n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, 
      n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, 
      n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, 
      n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, 
      n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, 
      n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, 
      n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, 
      n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, 
      n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, 
      n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, 
      n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, 
      n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, 
      n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, 
      n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, 
      n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, 
      n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, 
      n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, 
      n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, 
      n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, 
      n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, 
      n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, 
      n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, 
      n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, 
      n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, 
      n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, 
      n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, 
      n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, 
      n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, 
      n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, 
      n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, 
      n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, 
      n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, 
      n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, 
      n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, 
      n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, 
      n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, 
      n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, 
      n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, 
      n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, 
      n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, 
      n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, 
      n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, 
      n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, 
      n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, 
      n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, 
      n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, 
      n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, 
      n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, 
      n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, 
      n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, 
      n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, 
      n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, 
      n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, 
      n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, 
      n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, 
      n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, 
      n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, 
      n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, 
      n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, 
      n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, 
      n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, 
      n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, 
      n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, 
      n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, 
      n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, 
      n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, 
      n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, 
      n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, 
      n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, 
      n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, 
      n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, 
      n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, 
      n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, 
      n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, 
      n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, 
      n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, 
      n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, 
      n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, 
      n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, 
      n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, 
      n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, 
      n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, 
      n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, 
      n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, 
      n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, 
      n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, 
      n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, 
      n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, 
      n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, 
      n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, 
      n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, 
      n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, 
      n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, 
      n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, 
      n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, 
      n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, 
      n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, 
      n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, 
      n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, 
      n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, 
      n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, 
      n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, 
      n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, 
      n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, 
      n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, 
      n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, 
      n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, 
      n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, 
      n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, 
      n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, 
      n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, 
      n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, 
      n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, 
      n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, 
      n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, 
      n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, 
      n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, 
      n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, 
      n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, 
      n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, 
      n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, 
      n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, 
      n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, 
      n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, 
      n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, 
      n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, 
      n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, 
      n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, 
      n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, 
      n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, 
      n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, 
      n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, 
      n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, 
      n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, 
      n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, 
      n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, 
      n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, 
      n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, 
      n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, 
      n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, 
      n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, 
      n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, 
      n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, 
      n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, 
      n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, 
      n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, 
      n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, 
      n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, 
      n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, 
      n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, 
      n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, 
      n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, 
      n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, 
      n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, 
      n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, 
      n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, 
      n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, 
      n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, 
      n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, 
      n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, 
      n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, 
      n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, 
      n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, 
      n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, 
      n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, 
      n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, 
      n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, 
      n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, 
      n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, 
      n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, 
      n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, 
      n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, 
      n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, 
      n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, 
      n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, 
      n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, 
      n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, 
      n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, 
      n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, 
      n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, 
      n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, 
      n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, 
      n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, 
      n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, 
      n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, 
      n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, 
      n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, 
      n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, 
      n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, 
      n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, 
      n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, 
      n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, 
      n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, 
      n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, 
      n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, 
      n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, 
      n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, 
      n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, 
      n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, 
      n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, 
      n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, 
      n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, 
      n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, 
      n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, 
      n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, 
      n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, 
      n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, 
      n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, 
      n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, 
      n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, 
      n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, 
      n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, 
      n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, 
      n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, 
      n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, 
      n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, 
      n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, 
      n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, 
      n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, 
      n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, 
      n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, 
      n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, 
      n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, 
      n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, 
      n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, 
      n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, 
      n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, 
      n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, 
      n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, 
      n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, 
      n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, 
      n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, 
      n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, 
      n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, 
      n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, 
      n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, 
      n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, 
      n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, 
      n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, 
      n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, 
      n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, 
      n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, 
      n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, 
      n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, 
      n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, 
      n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, 
      n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, 
      n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, 
      n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, 
      n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, 
      n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, 
      n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, 
      n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, 
      n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, 
      n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, 
      n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, 
      n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, 
      n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, 
      n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, 
      n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, 
      n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, 
      n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, 
      n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, 
      n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, 
      n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, 
      n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, 
      n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, 
      n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, 
      n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, 
      n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, 
      n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, 
      n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, 
      n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, 
      n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, 
      n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, 
      n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, 
      n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, 
      n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, 
      n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, 
      n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, 
      n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, 
      n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, 
      n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, 
      n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, 
      n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, 
      n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, 
      n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, 
      n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, 
      n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, 
      n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, 
      n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, 
      n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, 
      n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, 
      n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, 
      n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, 
      n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, 
      n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, 
      n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, 
      n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, 
      n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, 
      n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, 
      n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, 
      n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, 
      n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, 
      n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, 
      n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, 
      n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, 
      n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, 
      n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, 
      n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, 
      n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, 
      n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, 
      n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, 
      n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, 
      n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, 
      n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, 
      n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, 
      n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, 
      n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, 
      n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, 
      n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, 
      n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, 
      n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, 
      n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, 
      n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, 
      n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, 
      n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, 
      n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, 
      n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, 
      n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, 
      n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, 
      n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, 
      n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, 
      n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, 
      n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, 
      n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, 
      n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, 
      n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, 
      n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, 
      n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, 
      n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, 
      n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, 
      n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, 
      n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, 
      n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, 
      n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, 
      n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, 
      n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, 
      n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, 
      n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, 
      n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, 
      n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, 
      n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, 
      n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, 
      n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, 
      n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, 
      n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, 
      n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, 
      n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, 
      n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, 
      n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, 
      n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, 
      n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, 
      n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, 
      n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, 
      n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, 
      n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, 
      n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, 
      n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, 
      n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, 
      n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, 
      n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, 
      n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, 
      n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, 
      n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, 
      n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, 
      n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, 
      n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, 
      n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, 
      n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, 
      n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, 
      n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, 
      n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, 
      n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, 
      n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, 
      n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, 
      n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, 
      n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, 
      n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, 
      n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, 
      n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, 
      n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, 
      n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, 
      n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, 
      n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, 
      n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, 
      n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, 
      n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, 
      n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, 
      n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, 
      n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, 
      n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, 
      n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, 
      n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, 
      n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, 
      n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, 
      n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, 
      n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, 
      n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, 
      n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, 
      n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, 
      n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, 
      n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, 
      n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, 
      n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, 
      n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, 
      n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, 
      n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, 
      n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, 
      n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, 
      n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, 
      n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, 
      n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, 
      n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, 
      n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, 
      n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, 
      n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, 
      n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, 
      n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, 
      n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, 
      n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, 
      n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, 
      n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, 
      n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, 
      n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, 
      n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, 
      n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, 
      n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, 
      n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, 
      n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, 
      n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, 
      n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, 
      n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, 
      n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, 
      n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, 
      n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, 
      n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, 
      n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, 
      n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, 
      n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, 
      n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, 
      n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, 
      n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, 
      n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, 
      n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, 
      n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, 
      n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, 
      n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, 
      n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, 
      n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, 
      n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, 
      n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, 
      n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, 
      n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, 
      n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, 
      n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, 
      n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, 
      n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, 
      n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, 
      n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, 
      n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, 
      n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, 
      n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, 
      n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, 
      n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, 
      n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, 
      n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, 
      n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, 
      n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, 
      n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, 
      n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, 
      n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, 
      n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, 
      n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, 
      n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, 
      n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, 
      n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, 
      n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, 
      n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, 
      n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, 
      n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, 
      n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, 
      n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, 
      n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, 
      n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, 
      n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, 
      n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618 : std_logic;

begin
   OUT1 <= ( OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, 
      OUT1_59_port, OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, 
      OUT1_54_port, OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, 
      OUT1_49_port, OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, 
      OUT1_44_port, OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, 
      OUT1_39_port, OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, 
      OUT1_34_port, OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, 
      OUT1_29_port, OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, 
      OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, 
      OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, 
      OUT1_14_port, OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, 
      OUT1_9_port, OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, 
      OUT1_4_port, OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port );
   MEM_BUS <= ( MEM_BUS_63_port, MEM_BUS_62_port, MEM_BUS_61_port, 
      MEM_BUS_60_port, MEM_BUS_59_port, MEM_BUS_58_port, MEM_BUS_57_port, 
      MEM_BUS_56_port, MEM_BUS_55_port, MEM_BUS_54_port, MEM_BUS_53_port, 
      MEM_BUS_52_port, MEM_BUS_51_port, MEM_BUS_50_port, MEM_BUS_49_port, 
      MEM_BUS_48_port, MEM_BUS_47_port, MEM_BUS_46_port, MEM_BUS_45_port, 
      MEM_BUS_44_port, MEM_BUS_43_port, MEM_BUS_42_port, MEM_BUS_41_port, 
      MEM_BUS_40_port, MEM_BUS_39_port, MEM_BUS_38_port, MEM_BUS_37_port, 
      MEM_BUS_36_port, MEM_BUS_35_port, MEM_BUS_34_port, MEM_BUS_33_port, 
      MEM_BUS_32_port, MEM_BUS_31_port, MEM_BUS_30_port, MEM_BUS_29_port, 
      MEM_BUS_28_port, MEM_BUS_27_port, MEM_BUS_26_port, MEM_BUS_25_port, 
      MEM_BUS_24_port, MEM_BUS_23_port, MEM_BUS_22_port, MEM_BUS_21_port, 
      MEM_BUS_20_port, MEM_BUS_19_port, MEM_BUS_18_port, MEM_BUS_17_port, 
      MEM_BUS_16_port, MEM_BUS_15_port, MEM_BUS_14_port, MEM_BUS_13_port, 
      MEM_BUS_12_port, MEM_BUS_11_port, MEM_BUS_10_port, MEM_BUS_9_port, 
      MEM_BUS_8_port, MEM_BUS_7_port, MEM_BUS_6_port, MEM_BUS_5_port, 
      MEM_BUS_4_port, MEM_BUS_3_port, MEM_BUS_2_port, MEM_BUS_1_port, 
      MEM_BUS_0_port );
   
   j_reg_0_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => n21416, QN => 
                           n5756);
   SWP_reg_31_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => n_1073, QN =>
                           n22794);
   SPILL_reg : DFF_X1 port map( D => n5643, CK => CLK, Q => SPILL, QN => n3236)
                           ;
   j_reg_31_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => n21455, QN => 
                           n5734);
   j_reg_30_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => n21453, QN => 
                           n5735);
   j_reg_29_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => n21449, QN => 
                           n5737);
   j_reg_28_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => n21446, QN => 
                           n5738);
   j_reg_27_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => n21442, QN => 
                           n5739);
   j_reg_26_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => n21441, QN => 
                           n5740);
   j_reg_25_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => n21439, QN => 
                           n5741);
   j_reg_24_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => n21437, QN => 
                           n5742);
   j_reg_23_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => n21434, QN => 
                           n5743);
   j_reg_22_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => n21433, QN => 
                           n5744);
   j_reg_21_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => n21436, QN => 
                           n5745);
   j_reg_20_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => n21435, QN => 
                           n5746);
   j_reg_19_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => n21030, QN => 
                           n5748);
   j_reg_18_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => n21430, QN => 
                           n5749);
   j_reg_17_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => n21431, QN => 
                           n5750);
   j_reg_16_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => n21432, QN => 
                           n_1074);
   j_reg_15_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => n21428, QN => 
                           n_1075);
   j_reg_14_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => n21029, QN => 
                           n5751);
   j_reg_13_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => n21426, QN => 
                           n5752);
   j_reg_12_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => n21427, QN => 
                           n5753);
   j_reg_11_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => n21028, QN => 
                           n5754);
   j_reg_10_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => n21425, QN => 
                           n_1076);
   j_reg_9_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => n21027, QN => 
                           n_1077);
   j_reg_8_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => n21424, QN => 
                           n5731);
   j_reg_7_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => n21423, QN => 
                           n_1078);
   j_reg_6_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => n21421, QN => 
                           n5732);
   j_reg_5_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => n21422, QN => 
                           n_1079);
   j_reg_4_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => n21420, QN => 
                           n5733);
   j_reg_3_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => n21418, QN => 
                           n5736);
   j_reg_2_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => n21419, QN => 
                           n5747);
   j_reg_1_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => n21417, QN => 
                           n5755);
   MEM_BUS_reg_0_inst : DFF_X1 port map( D => n22760, CK => CLK, Q => 
                           MEM_BUS_0_port, QN => n_1080);
   MEM_BUS_reg_6_inst : DFF_X1 port map( D => n22702, CK => CLK, Q => 
                           MEM_BUS_6_port, QN => n_1081);
   MEM_BUS_reg_5_inst : DFF_X1 port map( D => n22701, CK => CLK, Q => 
                           MEM_BUS_5_port, QN => n_1082);
   i_reg_0_inst : DFF_X1 port map( D => n13242, CK => CLK, Q => i_0_port, QN =>
                           n3242);
   i_reg_2_inst : DFF_X1 port map( D => n13240, CK => CLK, Q => i_2_port, QN =>
                           n3259);
   i_reg_3_inst : DFF_X1 port map( D => n13239, CK => CLK, Q => i_3_port, QN =>
                           n3253);
   i_reg_5_inst : DFF_X1 port map( D => n13237, CK => CLK, Q => i_5_port, QN =>
                           n3251);
   i_reg_6_inst : DFF_X1 port map( D => n13236, CK => CLK, Q => i_6_port, QN =>
                           n3258);
   i_reg_7_inst : DFF_X1 port map( D => n13235, CK => CLK, Q => i_7_port, QN =>
                           n3257);
   i_reg_10_inst : DFF_X1 port map( D => n13232, CK => CLK, Q => i_10_port, QN 
                           => n3241);
   i_reg_11_inst : DFF_X1 port map( D => n13231, CK => CLK, Q => i_11_port, QN 
                           => n3263);
   i_reg_12_inst : DFF_X1 port map( D => n13230, CK => CLK, Q => i_12_port, QN 
                           => n3262);
   i_reg_13_inst : DFF_X1 port map( D => n13229, CK => CLK, Q => i_13_port, QN 
                           => n3261);
   i_reg_14_inst : DFF_X1 port map( D => n13228, CK => CLK, Q => i_14_port, QN 
                           => n3260);
   i_reg_15_inst : DFF_X1 port map( D => n13227, CK => CLK, Q => i_15_port, QN 
                           => n3267);
   i_reg_16_inst : DFF_X1 port map( D => n13226, CK => CLK, Q => i_16_port, QN 
                           => n3266);
   i_reg_17_inst : DFF_X1 port map( D => n13225, CK => CLK, Q => i_17_port, QN 
                           => n3265);
   i_reg_18_inst : DFF_X1 port map( D => n13224, CK => CLK, Q => i_18_port, QN 
                           => n3264);
   i_reg_22_inst : DFF_X1 port map( D => n13220, CK => CLK, Q => i_22_port, QN 
                           => n3268);
   i_reg_23_inst : DFF_X1 port map( D => n13219, CK => CLK, Q => i_23_port, QN 
                           => n3246);
   i_reg_24_inst : DFF_X1 port map( D => n13218, CK => CLK, Q => i_24_port, QN 
                           => n3245);
   i_reg_25_inst : DFF_X1 port map( D => n13217, CK => CLK, Q => i_25_port, QN 
                           => n3244);
   i_reg_26_inst : DFF_X1 port map( D => n13216, CK => CLK, Q => i_26_port, QN 
                           => n3243);
   i_reg_27_inst : DFF_X1 port map( D => n13215, CK => CLK, Q => i_27_port, QN 
                           => n3250);
   i_reg_28_inst : DFF_X1 port map( D => n13214, CK => CLK, Q => i_28_port, QN 
                           => n3249);
   i_reg_29_inst : DFF_X1 port map( D => n13213, CK => CLK, Q => i_29_port, QN 
                           => n3248);
   i_reg_30_inst : DFF_X1 port map( D => n13212, CK => CLK, Q => i_30_port, QN 
                           => n3247);
   i_reg_31_inst : DFF_X1 port map( D => n13211, CK => CLK, Q => i_31_port, QN 
                           => n3254);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => OUT2(1), QN 
                           => n3141);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => OUT2(2), QN 
                           => n3140);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => OUT2(3), QN 
                           => n3139);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => OUT2(4), QN 
                           => n3138);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => OUT2(5), QN 
                           => n3137);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => OUT2(6), QN 
                           => n3136);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => OUT2(7), QN 
                           => n3135);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => OUT2(8), QN 
                           => n3134);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => OUT2(9), QN 
                           => n3133);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => OUT2(10), QN
                           => n3132);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => OUT2(11), QN
                           => n3131);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => OUT2(12), QN
                           => n3130);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => OUT2(13), QN
                           => n3129);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => OUT2(14), QN
                           => n3128);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => OUT2(15), QN
                           => n3127);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => OUT2(16), QN
                           => n3126);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => OUT2(17), QN
                           => n3125);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => OUT2(18), QN
                           => n3124);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => OUT2(19), QN
                           => n3123);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => OUT2(20), QN
                           => n3122);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => OUT2(21), QN
                           => n3121);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => OUT2(22), QN
                           => n3120);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => OUT2(23), QN
                           => n3119);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => OUT2(24), QN
                           => n3118);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => OUT2(25), QN
                           => n3117);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => OUT2(26), QN
                           => n3116);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => OUT2(27), QN
                           => n3115);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => OUT2(28), QN
                           => n3114);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => OUT2(29), QN
                           => n3113);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => OUT2(30), QN
                           => n3112);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => OUT2(31), QN
                           => n3111);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => OUT2(32), QN
                           => n3110);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => OUT2(33), QN
                           => n3109);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => OUT2(34), QN
                           => n3108);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => OUT2(35), QN
                           => n3107);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => OUT2(36), QN
                           => n3106);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => OUT2(37), QN
                           => n3105);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => OUT2(38), QN
                           => n3104);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => OUT2(39), QN
                           => n3103);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => OUT2(40), QN
                           => n3102);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => OUT2(41), QN
                           => n3101);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => OUT2(42), QN
                           => n3100);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => OUT2(43), QN
                           => n3099);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => OUT2(44), QN
                           => n3098);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => OUT2(45), QN
                           => n3097);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => OUT2(46), QN
                           => n3096);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => OUT2(47), QN
                           => n3095);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => OUT2(48), QN
                           => n3094);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => OUT2(49), QN
                           => n3093);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => OUT2(50), QN
                           => n3092);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => OUT2(51), QN
                           => n3091);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => OUT2(52), QN
                           => n3090);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => OUT2(53), QN
                           => n3089);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => OUT2(54), QN
                           => n3088);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => OUT2(55), QN
                           => n3087);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => OUT2(56), QN
                           => n3086);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => OUT2(57), QN
                           => n3085);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => OUT2(58), QN
                           => n3084);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => OUT2(59), QN
                           => n3083);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => OUT2(60), QN
                           => n3082);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => OUT2(61), QN
                           => n3081);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => OUT2(62), QN
                           => n3080);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => OUT2(63), QN
                           => n3079);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => OUT2(0), QN 
                           => n3078);
   FILL_reg : DFF_X1 port map( D => n5449, CK => CLK, Q => FILL, QN => n3077);
   SWP_reg_4_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => n_1083, QN => 
                           n22787);
   SWP_reg_6_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => n_1084, QN => 
                           n22791);
   SWP_reg_8_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => n_1085, QN => 
                           n22792);
   SWP_reg_14_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => n22534, QN =>
                           n22782);
   SWP_reg_20_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => n20750, QN =>
                           n22509);
   SWP_reg_21_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => n_1086, QN =>
                           n22786);
   SWP_reg_22_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => n_1087, QN =>
                           n22793);
   SWP_reg_23_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => n_1088, QN =>
                           n22795);
   SWP_reg_24_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => n_1089, QN =>
                           n22981);
   SWP_reg_25_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => n_1090, QN =>
                           n22783);
   SWP_reg_26_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => n_1091, QN =>
                           n22785);
   SWP_reg_27_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => n_1092, QN =>
                           n22789);
   SWP_reg_28_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => n_1093, QN =>
                           n22790);
   SWP_reg_9_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => n20732, QN => 
                           n22539);
   SWP_reg_7_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => n20734, QN => 
                           n22540);
   SWP_reg_5_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => n20736, QN => 
                           n22541);
   CWP_reg_1_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => CWP_1_port, QN
                           => n3044);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => 
                           n21750, QN => n18684);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => 
                           n21749, QN => n18685);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => 
                           n21709, QN => n18686);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => 
                           n21746, QN => n18687);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => 
                           n21745, QN => n18688);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => 
                           n21707, QN => n18689);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => 
                           n21742, QN => n18690);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => 
                           n21726, QN => n18691);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => 
                           n21705, QN => n18692);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => 
                           n21739, QN => n18693);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => 
                           n21738, QN => n18694);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => 
                           n21737, QN => n18695);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => 
                           n21702, QN => n18696);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => 
                           n21839, QN => n18697);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => 
                           n21701, QN => n18698);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => 
                           n21700, QN => n18699);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => 
                           n21724, QN => n18700);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => 
                           n21722, QN => n18701);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => 
                           n21721, QN => n18702);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => 
                           n21734, QN => n18703);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => 
                           n21720, QN => n18704);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => 
                           n21733, QN => n18705);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => 
                           n21697, QN => n18706);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => 
                           n21732, QN => n18707);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => 
                           n21835, QN => n18708);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => 
                           n21731, QN => n18709);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => 
                           n21714, QN => n18710);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => n21754
                           , QN => n18711);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => n21728
                           , QN => n18712);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => n21696
                           , QN => n18713);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => n21711
                           , QN => n18714);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => n21695
                           , QN => n18715);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => n21842
                           , QN => n18716);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => n21710
                           , QN => n18717);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => n21712
                           , QN => n18718);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => n21713
                           , QN => n18719);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => n21729
                           , QN => n18720);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => 
                           n21730, QN => n18721);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => 
                           n21715, QN => n18722);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => 
                           n21716, QN => n18723);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => 
                           n21717, QN => n18724);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => 
                           n21718, QN => n18725);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => 
                           n21719, QN => n18726);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => 
                           n21765, QN => n18727);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => 
                           n21698, QN => n18728);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => 
                           n21699, QN => n18729);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => 
                           n21735, QN => n18730);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => 
                           n21723, QN => n18731);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => 
                           n21837, QN => n18732);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => 
                           n21736, QN => n18733);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => 
                           n21838, QN => n18734);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => 
                           n21725, QN => n18735);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => 
                           n21836, QN => n18736);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => 
                           n21703, QN => n18737);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => 
                           n21704, QN => n18738);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => 
                           n21740, QN => n18739);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => 
                           n21741, QN => n18740);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => 
                           n21706, QN => n18741);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => 
                           n21743, QN => n18742);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => 
                           n21744, QN => n18743);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => 
                           n21708, QN => n18744);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => 
                           n21747, QN => n18745);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => 
                           n21748, QN => n18746);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => 
                           n21727, QN => n18747);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => 
                           n21694, QN => n18748);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => 
                           n21693, QN => n18749);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => 
                           n21653, QN => n18750);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => 
                           n21690, QN => n18751);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => 
                           n21689, QN => n18752);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => 
                           n21651, QN => n18753);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => 
                           n21686, QN => n18754);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => 
                           n21670, QN => n18755);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => 
                           n21649, QN => n18756);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => 
                           n21683, QN => n18757);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => 
                           n21682, QN => n18758);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => 
                           n21681, QN => n18759);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => 
                           n21646, QN => n18760);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => 
                           n21834, QN => n18761);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => 
                           n21645, QN => n18762);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => 
                           n21644, QN => n18763);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => 
                           n21668, QN => n18764);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => 
                           n21666, QN => n18765);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => 
                           n21665, QN => n18766);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => 
                           n21678, QN => n18767);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => 
                           n21664, QN => n18768);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => 
                           n21677, QN => n18769);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => 
                           n21642, QN => n18770);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => 
                           n21676, QN => n18771);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => 
                           n21830, QN => n18772);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => 
                           n21675, QN => n18773);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => 
                           n21658, QN => n18774);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => n21751
                           , QN => n18775);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => n21672
                           , QN => n18776);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => n21641
                           , QN => n18777);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => n21655
                           , QN => n18778);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => n21640
                           , QN => n18779);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => n21843
                           , QN => n18780);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => n21654
                           , QN => n18781);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => n21656
                           , QN => n18782);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => n21657
                           , QN => n18783);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => n21673
                           , QN => n18784);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => 
                           n21674, QN => n18785);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => 
                           n21659, QN => n18786);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => 
                           n21660, QN => n18787);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n5310, CK => CLK, Q => 
                           n21661, QN => n18788);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n5309, CK => CLK, Q => 
                           n21662, QN => n18789);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n5308, CK => CLK, Q => 
                           n21663, QN => n18790);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n5307, CK => CLK, Q => 
                           n21764, QN => n18791);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n5306, CK => CLK, Q => 
                           n21639, QN => n18792);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n5305, CK => CLK, Q => 
                           n21643, QN => n18793);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n5304, CK => CLK, Q => 
                           n21679, QN => n18794);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n5303, CK => CLK, Q => 
                           n21667, QN => n18795);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n5302, CK => CLK, Q => 
                           n21832, QN => n18796);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n5301, CK => CLK, Q => 
                           n21680, QN => n18797);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n5300, CK => CLK, Q => 
                           n21833, QN => n18798);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n5299, CK => CLK, Q => 
                           n21669, QN => n18799);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n5298, CK => CLK, Q => 
                           n21831, QN => n18800);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n5297, CK => CLK, Q => 
                           n21647, QN => n18801);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n5296, CK => CLK, Q => 
                           n21648, QN => n18802);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n5295, CK => CLK, Q => 
                           n21684, QN => n18803);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n5294, CK => CLK, Q => 
                           n21685, QN => n18804);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n5293, CK => CLK, Q => 
                           n21650, QN => n18805);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n5292, CK => CLK, Q => 
                           n21687, QN => n18806);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n5291, CK => CLK, Q => 
                           n21688, QN => n18807);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n5290, CK => CLK, Q => 
                           n21652, QN => n18808);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n5289, CK => CLK, Q => 
                           n21691, QN => n18809);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n5288, CK => CLK, Q => 
                           n21692, QN => n18810);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n5287, CK => CLK, Q => 
                           n21671, QN => n18811);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n5286, CK => CLK, Q => 
                           n21265, QN => n18812);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n5285, CK => CLK, Q => 
                           n21264, QN => n18813);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n5284, CK => CLK, Q => 
                           n21224, QN => n18814);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n5283, CK => CLK, Q => 
                           n21261, QN => n18815);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n5282, CK => CLK, Q => 
                           n21243, QN => n18816);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n5281, CK => CLK, Q => 
                           n21222, QN => n18817);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n5280, CK => CLK, Q => 
                           n21258, QN => n18818);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n5279, CK => CLK, Q => 
                           n21241, QN => n18819);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n5278, CK => CLK, Q => 
                           n21220, QN => n18820);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n5277, CK => CLK, Q => 
                           n21255, QN => n18821);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n5276, CK => CLK, Q => 
                           n21254, QN => n18822);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n5275, CK => CLK, Q => 
                           n21253, QN => n18823);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n5274, CK => CLK, Q => 
                           n21217, QN => n18824);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n5273, CK => CLK, Q => 
                           n21283, QN => n18825);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n5272, CK => CLK, Q => 
                           n21216, QN => n18826);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n5271, CK => CLK, Q => 
                           n21215, QN => n18827);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n5270, CK => CLK, Q => 
                           n21239, QN => n18828);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n5269, CK => CLK, Q => 
                           n21237, QN => n18829);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n5268, CK => CLK, Q => 
                           n21236, QN => n18830);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n5267, CK => CLK, Q => 
                           n21250, QN => n18831);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n5266, CK => CLK, Q => 
                           n21235, QN => n18832);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n5265, CK => CLK, Q => 
                           n21249, QN => n18833);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n5264, CK => CLK, Q => 
                           n21212, QN => n18834);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n5263, CK => CLK, Q => 
                           n21248, QN => n18835);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n5262, CK => CLK, Q => 
                           n21279, QN => n18836);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n5261, CK => CLK, Q => 
                           n21247, QN => n18837);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n5260, CK => CLK, Q => 
                           n21229, QN => n18838);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n5259, CK => CLK, Q => n21266
                           , QN => n18839);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n5258, CK => CLK, Q => n21244
                           , QN => n18840);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n5257, CK => CLK, Q => n21211
                           , QN => n18841);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n5256, CK => CLK, Q => n21226
                           , QN => n18842);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n5255, CK => CLK, Q => n21210
                           , QN => n18843);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n5254, CK => CLK, Q => n21285
                           , QN => n18844);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n5253, CK => CLK, Q => n21225
                           , QN => n18845);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n5252, CK => CLK, Q => n21227
                           , QN => n18846);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n5251, CK => CLK, Q => n21228
                           , QN => n18847);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n5250, CK => CLK, Q => n21245
                           , QN => n18848);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n5249, CK => CLK, Q => 
                           n21246, QN => n18849);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n5248, CK => CLK, Q => 
                           n21230, QN => n18850);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n5247, CK => CLK, Q => 
                           n21231, QN => n18851);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n5246, CK => CLK, Q => 
                           n21232, QN => n18852);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n5245, CK => CLK, Q => 
                           n21233, QN => n18853);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n5244, CK => CLK, Q => 
                           n21234, QN => n18854);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n5243, CK => CLK, Q => 
                           n21274, QN => n18855);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n5242, CK => CLK, Q => 
                           n21213, QN => n18856);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n5241, CK => CLK, Q => 
                           n21214, QN => n18857);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n5240, CK => CLK, Q => 
                           n21251, QN => n18858);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n5239, CK => CLK, Q => 
                           n21238, QN => n18859);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n5238, CK => CLK, Q => 
                           n21281, QN => n18860);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n5237, CK => CLK, Q => 
                           n21252, QN => n18861);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n5236, CK => CLK, Q => 
                           n21282, QN => n18862);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n5235, CK => CLK, Q => 
                           n21240, QN => n18863);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n5234, CK => CLK, Q => 
                           n21280, QN => n18864);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n5233, CK => CLK, Q => 
                           n21218, QN => n18865);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n5232, CK => CLK, Q => 
                           n21219, QN => n18866);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n5231, CK => CLK, Q => 
                           n21256, QN => n18867);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n5230, CK => CLK, Q => 
                           n21257, QN => n18868);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n5229, CK => CLK, Q => 
                           n21221, QN => n18869);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n5228, CK => CLK, Q => 
                           n21259, QN => n18870);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n5227, CK => CLK, Q => 
                           n21260, QN => n18871);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n5226, CK => CLK, Q => 
                           n21223, QN => n18872);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n5225, CK => CLK, Q => 
                           n21262, QN => n18873);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n5224, CK => CLK, Q => 
                           n21263, QN => n18874);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n5223, CK => CLK, Q => 
                           n21242, QN => n18875);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n5222, CK => CLK, Q => 
                           n20954, QN => n18876);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n5221, CK => CLK, Q => 
                           n20953, QN => n18877);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n5220, CK => CLK, Q => 
                           n20913, QN => n18878);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n5219, CK => CLK, Q => 
                           n20950, QN => n18879);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n5218, CK => CLK, Q => 
                           n20949, QN => n18880);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n5217, CK => CLK, Q => 
                           n20911, QN => n18881);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n5216, CK => CLK, Q => 
                           n20946, QN => n18882);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n5215, CK => CLK, Q => 
                           n20930, QN => n18883);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n5214, CK => CLK, Q => 
                           n20909, QN => n18884);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n5213, CK => CLK, Q => 
                           n20943, QN => n18885);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n5212, CK => CLK, Q => 
                           n20942, QN => n18886);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n5211, CK => CLK, Q => 
                           n20941, QN => n18887);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n5210, CK => CLK, Q => 
                           n20906, QN => n18888);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n5209, CK => CLK, Q => 
                           n20961, QN => n18889);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n5208, CK => CLK, Q => 
                           n20905, QN => n18890);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n5207, CK => CLK, Q => 
                           n20904, QN => n18891);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n5206, CK => CLK, Q => 
                           n20928, QN => n18892);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n5205, CK => CLK, Q => 
                           n20926, QN => n18893);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n5204, CK => CLK, Q => 
                           n20925, QN => n18894);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n5203, CK => CLK, Q => 
                           n20938, QN => n18895);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n5202, CK => CLK, Q => 
                           n20924, QN => n18896);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n5201, CK => CLK, Q => 
                           n20937, QN => n18897);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n5200, CK => CLK, Q => 
                           n20902, QN => n18898);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n5199, CK => CLK, Q => 
                           n20936, QN => n18899);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n5198, CK => CLK, Q => 
                           n20957, QN => n18900);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n5197, CK => CLK, Q => 
                           n20935, QN => n18901);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n5196, CK => CLK, Q => 
                           n20918, QN => n18902);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n5195, CK => CLK, Q => n20955
                           , QN => n18903);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n5194, CK => CLK, Q => n20932
                           , QN => n18904);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n5193, CK => CLK, Q => n20901
                           , QN => n18905);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n5192, CK => CLK, Q => n20915
                           , QN => n18906);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n5191, CK => CLK, Q => n20900
                           , QN => n18907);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n5190, CK => CLK, Q => n20962
                           , QN => n18908);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n5189, CK => CLK, Q => n20914
                           , QN => n18909);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n5188, CK => CLK, Q => n20916
                           , QN => n18910);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n5187, CK => CLK, Q => n20917
                           , QN => n18911);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n5186, CK => CLK, Q => n20933
                           , QN => n18912);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n5185, CK => CLK, Q => 
                           n20934, QN => n18913);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n5184, CK => CLK, Q => 
                           n20919, QN => n18914);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n5183, CK => CLK, Q => 
                           n20920, QN => n18915);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n5182, CK => CLK, Q => 
                           n20921, QN => n18916);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n5181, CK => CLK, Q => 
                           n20922, QN => n18917);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n5180, CK => CLK, Q => 
                           n20923, QN => n18918);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n5179, CK => CLK, Q => 
                           n20956, QN => n18919);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n5178, CK => CLK, Q => 
                           n20899, QN => n18920);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n5177, CK => CLK, Q => 
                           n20903, QN => n18921);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n5176, CK => CLK, Q => 
                           n20939, QN => n18922);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n5175, CK => CLK, Q => 
                           n20927, QN => n18923);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n5174, CK => CLK, Q => 
                           n20959, QN => n18924);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n5173, CK => CLK, Q => 
                           n20940, QN => n18925);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n5172, CK => CLK, Q => 
                           n20960, QN => n18926);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n5171, CK => CLK, Q => 
                           n20929, QN => n18927);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n5170, CK => CLK, Q => 
                           n20958, QN => n18928);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n5169, CK => CLK, Q => 
                           n20907, QN => n18929);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n5168, CK => CLK, Q => 
                           n20908, QN => n18930);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n5167, CK => CLK, Q => 
                           n20944, QN => n18931);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n5166, CK => CLK, Q => 
                           n20945, QN => n18932);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n5165, CK => CLK, Q => 
                           n20910, QN => n18933);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n5164, CK => CLK, Q => 
                           n20947, QN => n18934);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n5163, CK => CLK, Q => 
                           n20948, QN => n18935);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n5162, CK => CLK, Q => 
                           n20912, QN => n18936);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n5161, CK => CLK, Q => 
                           n20951, QN => n18937);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n5160, CK => CLK, Q => 
                           n20952, QN => n18938);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n5159, CK => CLK, Q => 
                           n20931, QN => n18939);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n5158, CK => CLK, Q => 
                           n22229, QN => n18940);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n5157, CK => CLK, Q => 
                           n22230, QN => n18941);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n5156, CK => CLK, Q => 
                           n22231, QN => n18942);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n5155, CK => CLK, Q => 
                           n22232, QN => n18943);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n5154, CK => CLK, Q => 
                           n22233, QN => n18944);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n5153, CK => CLK, Q => 
                           n22234, QN => n18945);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n5152, CK => CLK, Q => 
                           n22227, QN => n18946);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n5151, CK => CLK, Q => 
                           n22235, QN => n18947);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n5150, CK => CLK, Q => 
                           n22236, QN => n18948);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n5149, CK => CLK, Q => 
                           n22237, QN => n18949);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n5148, CK => CLK, Q => 
                           n22238, QN => n18950);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n5147, CK => CLK, Q => 
                           n22239, QN => n18951);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n5146, CK => CLK, Q => 
                           n22240, QN => n18952);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n5145, CK => CLK, Q => 
                           n22241, QN => n18953);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n5144, CK => CLK, Q => 
                           n22242, QN => n18954);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n5143, CK => CLK, Q => 
                           n22243, QN => n18955);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n5142, CK => CLK, Q => 
                           n22244, QN => n18956);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n5141, CK => CLK, Q => 
                           n22245, QN => n18957);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n5140, CK => CLK, Q => 
                           n22228, QN => n18958);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n5139, CK => CLK, Q => 
                           n22246, QN => n18959);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n5138, CK => CLK, Q => 
                           n22247, QN => n18960);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n5137, CK => CLK, Q => 
                           n22248, QN => n18961);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n5136, CK => CLK, Q => 
                           n22249, QN => n18962);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n5135, CK => CLK, Q => 
                           n22261, QN => n18963);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n5134, CK => CLK, Q => 
                           n22250, QN => n18964);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n5133, CK => CLK, Q => 
                           n22251, QN => n18965);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n5132, CK => CLK, Q => 
                           n22252, QN => n18966);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n5131, CK => CLK, Q => n22253
                           , QN => n18967);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n5130, CK => CLK, Q => n22254
                           , QN => n18968);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n5129, CK => CLK, Q => n22262
                           , QN => n18969);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n5128, CK => CLK, Q => n22255
                           , QN => n18970);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n5127, CK => CLK, Q => n22256
                           , QN => n18971);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n5126, CK => CLK, Q => n22226
                           , QN => n18972);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n5125, CK => CLK, Q => n22257
                           , QN => n18973);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n5124, CK => CLK, Q => n22258
                           , QN => n18974);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n5123, CK => CLK, Q => n22263
                           , QN => n18975);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n5122, CK => CLK, Q => n22264
                           , QN => n18976);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n5121, CK => CLK, Q => 
                           n22265, QN => n18977);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n5120, CK => CLK, Q => 
                           n22266, QN => n18978);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n5119, CK => CLK, Q => 
                           n22267, QN => n18979);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n5118, CK => CLK, Q => 
                           n22268, QN => n18980);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n5117, CK => CLK, Q => 
                           n22259, QN => n18981);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n5116, CK => CLK, Q => 
                           n22269, QN => n18982);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n5115, CK => CLK, Q => 
                           n22270, QN => n18983);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n5114, CK => CLK, Q => 
                           n22271, QN => n18984);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n5113, CK => CLK, Q => 
                           n22272, QN => n18985);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n5112, CK => CLK, Q => 
                           n22273, QN => n18986);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n5111, CK => CLK, Q => 
                           n22274, QN => n18987);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n5110, CK => CLK, Q => 
                           n22275, QN => n18988);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n5109, CK => CLK, Q => 
                           n22276, QN => n18989);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n5108, CK => CLK, Q => 
                           n22277, QN => n18990);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n5107, CK => CLK, Q => 
                           n22278, QN => n18991);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n5106, CK => CLK, Q => 
                           n22279, QN => n18992);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n5105, CK => CLK, Q => 
                           n22260, QN => n18993);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n5104, CK => CLK, Q => 
                           n22280, QN => n18994);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n5103, CK => CLK, Q => 
                           n22281, QN => n18995);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n5102, CK => CLK, Q => 
                           n22282, QN => n18996);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n5101, CK => CLK, Q => 
                           n22283, QN => n18997);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n5100, CK => CLK, Q => 
                           n22284, QN => n18998);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n5099, CK => CLK, Q => 
                           n22285, QN => n18999);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n5098, CK => CLK, Q => 
                           n22286, QN => n19000);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n5097, CK => CLK, Q => 
                           n22287, QN => n19001);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n5096, CK => CLK, Q => 
                           n22288, QN => n19002);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n5095, CK => CLK, Q => 
                           n22289, QN => n19003);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n5094, CK => CLK, Q => 
                           n22057, QN => n19004);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n5093, CK => CLK, Q => 
                           n22182, QN => n19005);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n5092, CK => CLK, Q => 
                           n22056, QN => n19006);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n5091, CK => CLK, Q => 
                           n22179, QN => n19007);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n5090, CK => CLK, Q => 
                           n22036, QN => n19008);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n5089, CK => CLK, Q => 
                           n22055, QN => n19009);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n5088, CK => CLK, Q => 
                           n22175, QN => n19010);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n5087, CK => CLK, Q => 
                           n22173, QN => n19011);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n5086, CK => CLK, Q => 
                           n22172, QN => n19012);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n5085, CK => CLK, Q => 
                           n22170, QN => n19013);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n5084, CK => CLK, Q => 
                           n22168, QN => n19014);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n5083, CK => CLK, Q => 
                           n22053, QN => n19015);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n5082, CK => CLK, Q => 
                           n22165, QN => n19016);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n5081, CK => CLK, Q => 
                           n22164, QN => n19017);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n5080, CK => CLK, Q => 
                           n22162, QN => n19018);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n5079, CK => CLK, Q => 
                           n22051, QN => n19019);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n5078, CK => CLK, Q => 
                           n22049, QN => n19020);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n5077, CK => CLK, Q => 
                           n22047, QN => n19021);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n5076, CK => CLK, Q => 
                           n22045, QN => n19022);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n5075, CK => CLK, Q => 
                           n22043, QN => n19023);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n5074, CK => CLK, Q => 
                           n22159, QN => n19024);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n5073, CK => CLK, Q => 
                           n22158, QN => n19025);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n5072, CK => CLK, Q => 
                           n22156, QN => n19026);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n5071, CK => CLK, Q => 
                           n22155, QN => n19027);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n5070, CK => CLK, Q => 
                           n22040, QN => n19028);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n5069, CK => CLK, Q => 
                           n22152, QN => n19029);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n5068, CK => CLK, Q => 
                           n22150, QN => n19030);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n5067, CK => CLK, Q => n22039
                           , QN => n19031);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n5066, CK => CLK, Q => n22147
                           , QN => n19032);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n5065, CK => CLK, Q => n22145
                           , QN => n19033);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n5064, CK => CLK, Q => n22038
                           , QN => n19034);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n5063, CK => CLK, Q => n22143
                           , QN => n19035);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n5062, CK => CLK, Q => n22291
                           , QN => n19036);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n5061, CK => CLK, Q => n22037
                           , QN => n19037);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n5060, CK => CLK, Q => n22144
                           , QN => n19038);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n5059, CK => CLK, Q => n22146
                           , QN => n19039);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n5058, CK => CLK, Q => n22148
                           , QN => n19040);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n5057, CK => CLK, Q => 
                           n22149, QN => n19041);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n5056, CK => CLK, Q => 
                           n22151, QN => n19042);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n5055, CK => CLK, Q => 
                           n22153, QN => n19043);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n5054, CK => CLK, Q => 
                           n22154, QN => n19044);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n5053, CK => CLK, Q => 
                           n22041, QN => n19045);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n5052, CK => CLK, Q => 
                           n22157, QN => n19046);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n5051, CK => CLK, Q => 
                           n22042, QN => n19047);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n5050, CK => CLK, Q => 
                           n22160, QN => n19048);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n5049, CK => CLK, Q => 
                           n22044, QN => n19049);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n5048, CK => CLK, Q => 
                           n22046, QN => n19050);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n5047, CK => CLK, Q => 
                           n22048, QN => n19051);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n5046, CK => CLK, Q => 
                           n22050, QN => n19052);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n5045, CK => CLK, Q => 
                           n22161, QN => n19053);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n5044, CK => CLK, Q => 
                           n22163, QN => n19054);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n5043, CK => CLK, Q => 
                           n22052, QN => n19055);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n5042, CK => CLK, Q => 
                           n22166, QN => n19056);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n5041, CK => CLK, Q => 
                           n22167, QN => n19057);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n5040, CK => CLK, Q => 
                           n22169, QN => n19058);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n5039, CK => CLK, Q => 
                           n22171, QN => n19059);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n5038, CK => CLK, Q => 
                           n22054, QN => n19060);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n5037, CK => CLK, Q => 
                           n22174, QN => n19061);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n5036, CK => CLK, Q => 
                           n22176, QN => n19062);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n5035, CK => CLK, Q => 
                           n22177, QN => n19063);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n5034, CK => CLK, Q => 
                           n22178, QN => n19064);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n5033, CK => CLK, Q => 
                           n22180, QN => n19065);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n5032, CK => CLK, Q => 
                           n22181, QN => n19066);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n5031, CK => CLK, Q => 
                           n22183, QN => n19067);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n5030, CK => CLK, Q => 
                           n22481, QN => n19068);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n5029, CK => CLK, Q => 
                           n22479, QN => n19069);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n5028, CK => CLK, Q => 
                           n22477, QN => n19070);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n5027, CK => CLK, Q => 
                           n22475, QN => n19071);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n5026, CK => CLK, Q => 
                           n22451, QN => n19072);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n5025, CK => CLK, Q => 
                           n22450, QN => n19073);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n5024, CK => CLK, Q => 
                           n22449, QN => n19074);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n5023, CK => CLK, Q => 
                           n22447, QN => n19075);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n5022, CK => CLK, Q => 
                           n22445, QN => n19076);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n5021, CK => CLK, Q => 
                           n22443, QN => n19077);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n5020, CK => CLK, Q => 
                           n22441, QN => n19078);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n5019, CK => CLK, Q => 
                           n22471, QN => n19079);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n5018, CK => CLK, Q => 
                           n22470, QN => n19080);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n5017, CK => CLK, Q => 
                           n22469, QN => n19081);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n5016, CK => CLK, Q => 
                           n22467, QN => n19082);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n5015, CK => CLK, Q => 
                           n22465, QN => n19083);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n5014, CK => CLK, Q => 
                           n22437, QN => n19084);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n5013, CK => CLK, Q => 
                           n22436, QN => n19085);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n5012, CK => CLK, Q => 
                           n22435, QN => n19086);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n5011, CK => CLK, Q => 
                           n22433, QN => n19087);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n5010, CK => CLK, Q => 
                           n22431, QN => n19088);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n5009, CK => CLK, Q => 
                           n22429, QN => n19089);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n5008, CK => CLK, Q => 
                           n22427, QN => n19090);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n5007, CK => CLK, Q => 
                           n22461, QN => n19091);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n5006, CK => CLK, Q => 
                           n22460, QN => n19092);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n5005, CK => CLK, Q => 
                           n22459, QN => n19093);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n5004, CK => CLK, Q => 
                           n22457, QN => n19094);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n5003, CK => CLK, Q => n22455
                           , QN => n19095);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n5002, CK => CLK, Q => n22423
                           , QN => n19096);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n5001, CK => CLK, Q => n22422
                           , QN => n19097);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n5000, CK => CLK, Q => n22420
                           , QN => n19098);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n4999, CK => CLK, Q => n22418
                           , QN => n19099);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n4998, CK => CLK, Q => n22452
                           , QN => n19100);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n4997, CK => CLK, Q => n22419
                           , QN => n19101);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n4996, CK => CLK, Q => n22421
                           , QN => n19102);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n4995, CK => CLK, Q => n22453
                           , QN => n19103);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n4994, CK => CLK, Q => n22454
                           , QN => n19104);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n4993, CK => CLK, Q => 
                           n22456, QN => n19105);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n4992, CK => CLK, Q => 
                           n22458, QN => n19106);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n4991, CK => CLK, Q => 
                           n22424, QN => n19107);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n4990, CK => CLK, Q => 
                           n22425, QN => n19108);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n4989, CK => CLK, Q => 
                           n22426, QN => n19109);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n4988, CK => CLK, Q => 
                           n22428, QN => n19110);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n4987, CK => CLK, Q => 
                           n22430, QN => n19111);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n4986, CK => CLK, Q => 
                           n22432, QN => n19112);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n4985, CK => CLK, Q => 
                           n22434, QN => n19113);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n4984, CK => CLK, Q => 
                           n22462, QN => n19114);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n4983, CK => CLK, Q => 
                           n22463, QN => n19115);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n4982, CK => CLK, Q => 
                           n22464, QN => n19116);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n4981, CK => CLK, Q => 
                           n22466, QN => n19117);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n4980, CK => CLK, Q => 
                           n22468, QN => n19118);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n4979, CK => CLK, Q => 
                           n22438, QN => n19119);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n4978, CK => CLK, Q => 
                           n22439, QN => n19120);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n4977, CK => CLK, Q => 
                           n22440, QN => n19121);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n4976, CK => CLK, Q => 
                           n22442, QN => n19122);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n4975, CK => CLK, Q => 
                           n22444, QN => n19123);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n4974, CK => CLK, Q => 
                           n22446, QN => n19124);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n4973, CK => CLK, Q => 
                           n22448, QN => n19125);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n4972, CK => CLK, Q => 
                           n22472, QN => n19126);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n4971, CK => CLK, Q => 
                           n22473, QN => n19127);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n4970, CK => CLK, Q => 
                           n22474, QN => n19128);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n4969, CK => CLK, Q => 
                           n22476, QN => n19129);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n4968, CK => CLK, Q => 
                           n22478, QN => n19130);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n4967, CK => CLK, Q => 
                           n22480, QN => n19131);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n4966, CK => CLK, Q => 
                           n21825, QN => n19132);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n4965, CK => CLK, Q => 
                           n21823, QN => n19133);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n4964, CK => CLK, Q => 
                           n21821, QN => n19134);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n4963, CK => CLK, Q => 
                           n21819, QN => n19135);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n4962, CK => CLK, Q => 
                           n21817, QN => n19136);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n4961, CK => CLK, Q => 
                           n21815, QN => n19137);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n4960, CK => CLK, Q => 
                           n21813, QN => n19138);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n4959, CK => CLK, Q => 
                           n21811, QN => n19139);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n4958, CK => CLK, Q => 
                           n21809, QN => n19140);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n4957, CK => CLK, Q => 
                           n21807, QN => n19141);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n4956, CK => CLK, Q => 
                           n21805, QN => n19142);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n4955, CK => CLK, Q => 
                           n21803, QN => n19143);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n4954, CK => CLK, Q => 
                           n21801, QN => n19144);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n4953, CK => CLK, Q => 
                           n21799, QN => n19145);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n4952, CK => CLK, Q => 
                           n21797, QN => n19146);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n4951, CK => CLK, Q => 
                           n21795, QN => n19147);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n4950, CK => CLK, Q => 
                           n21793, QN => n19148);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n4949, CK => CLK, Q => 
                           n21791, QN => n19149);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n4948, CK => CLK, Q => 
                           n21789, QN => n19150);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n4947, CK => CLK, Q => 
                           n21787, QN => n19151);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n4946, CK => CLK, Q => 
                           n21785, QN => n19152);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n4945, CK => CLK, Q => 
                           n21783, QN => n19153);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n4944, CK => CLK, Q => 
                           n21781, QN => n19154);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n4943, CK => CLK, Q => 
                           n21779, QN => n19155);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n4942, CK => CLK, Q => 
                           n21777, QN => n19156);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n4941, CK => CLK, Q => 
                           n21775, QN => n19157);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n4940, CK => CLK, Q => 
                           n21773, QN => n19158);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n4939, CK => CLK, Q => n21771
                           , QN => n19159);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n4938, CK => CLK, Q => n21769
                           , QN => n19160);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n4937, CK => CLK, Q => n21767
                           , QN => n19161);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n4936, CK => CLK, Q => n21828
                           , QN => n19162);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n4935, CK => CLK, Q => n21826
                           , QN => n19163);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n4934, CK => CLK, Q => n21766
                           , QN => n19164);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n4933, CK => CLK, Q => n21827
                           , QN => n19165);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n4932, CK => CLK, Q => n21829
                           , QN => n19166);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n4931, CK => CLK, Q => n21768
                           , QN => n19167);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n4930, CK => CLK, Q => n21770
                           , QN => n19168);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n4929, CK => CLK, Q => 
                           n21772, QN => n19169);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n4928, CK => CLK, Q => 
                           n21774, QN => n19170);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n4927, CK => CLK, Q => 
                           n21776, QN => n19171);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n4926, CK => CLK, Q => 
                           n21778, QN => n19172);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n4925, CK => CLK, Q => 
                           n21780, QN => n19173);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n4924, CK => CLK, Q => 
                           n21782, QN => n19174);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n4923, CK => CLK, Q => 
                           n21784, QN => n19175);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n4922, CK => CLK, Q => 
                           n21786, QN => n19176);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n4921, CK => CLK, Q => 
                           n21788, QN => n19177);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n4920, CK => CLK, Q => 
                           n21790, QN => n19178);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n4919, CK => CLK, Q => 
                           n21792, QN => n19179);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n4918, CK => CLK, Q => 
                           n21794, QN => n19180);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n4917, CK => CLK, Q => 
                           n21796, QN => n19181);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n4916, CK => CLK, Q => 
                           n21798, QN => n19182);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n4915, CK => CLK, Q => 
                           n21800, QN => n19183);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n4914, CK => CLK, Q => 
                           n21802, QN => n19184);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n4913, CK => CLK, Q => 
                           n21804, QN => n19185);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n4912, CK => CLK, Q => 
                           n21806, QN => n19186);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n4911, CK => CLK, Q => 
                           n21808, QN => n19187);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n4910, CK => CLK, Q => 
                           n21810, QN => n19188);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n4909, CK => CLK, Q => 
                           n21812, QN => n19189);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n4908, CK => CLK, Q => 
                           n21814, QN => n19190);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n4907, CK => CLK, Q => 
                           n21816, QN => n19191);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n4906, CK => CLK, Q => 
                           n21818, QN => n19192);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n4905, CK => CLK, Q => 
                           n21820, QN => n19193);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n4904, CK => CLK, Q => 
                           n21822, QN => n19194);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n4903, CK => CLK, Q => 
                           n21824, QN => n19195);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n4902, CK => CLK, Q => 
                           n21635, QN => n19196);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n4901, CK => CLK, Q => 
                           n21634, QN => n19197);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n4900, CK => CLK, Q => 
                           n21593, QN => n19198);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n4899, CK => CLK, Q => 
                           n21629, QN => n19199);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n4898, CK => CLK, Q => 
                           n21628, QN => n19200);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n4897, CK => CLK, Q => 
                           n21591, QN => n19201);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n4896, CK => CLK, Q => 
                           n21625, QN => n19202);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n4895, CK => CLK, Q => 
                           n21610, QN => n19203);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n4894, CK => CLK, Q => 
                           n21589, QN => n19204);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n4893, CK => CLK, Q => 
                           n21622, QN => n19205);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n4892, CK => CLK, Q => 
                           n21621, QN => n19206);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n4891, CK => CLK, Q => 
                           n21620, QN => n19207);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n4890, CK => CLK, Q => 
                           n21586, QN => n19208);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n4889, CK => CLK, Q => 
                           n21762, QN => n19209);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n4888, CK => CLK, Q => 
                           n21585, QN => n19210);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n4887, CK => CLK, Q => 
                           n21584, QN => n19211);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n4886, CK => CLK, Q => 
                           n21608, QN => n19212);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n4885, CK => CLK, Q => 
                           n21606, QN => n19213);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n4884, CK => CLK, Q => 
                           n21605, QN => n19214);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n4883, CK => CLK, Q => 
                           n21617, QN => n19215);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n4882, CK => CLK, Q => 
                           n21604, QN => n19216);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n4881, CK => CLK, Q => 
                           n21616, QN => n19217);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n4880, CK => CLK, Q => 
                           n21581, QN => n19218);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n4879, CK => CLK, Q => 
                           n21615, QN => n19219);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n4878, CK => CLK, Q => 
                           n21758, QN => n19220);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n4877, CK => CLK, Q => 
                           n21614, QN => n19221);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n4876, CK => CLK, Q => 
                           n21598, QN => n19222);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n4875, CK => CLK, Q => n21636
                           , QN => n19223);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n4874, CK => CLK, Q => n21611
                           , QN => n19224);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n4873, CK => CLK, Q => n21580
                           , QN => n19225);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n4872, CK => CLK, Q => n21595
                           , QN => n19226);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n4871, CK => CLK, Q => n21579
                           , QN => n19227);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n4870, CK => CLK, Q => n21840
                           , QN => n19228);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n4869, CK => CLK, Q => n21594
                           , QN => n19229);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n4868, CK => CLK, Q => n21596
                           , QN => n19230);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n4867, CK => CLK, Q => n21597
                           , QN => n19231);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n4866, CK => CLK, Q => n21612
                           , QN => n19232);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n4865, CK => CLK, Q => 
                           n21613, QN => n19233);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n4864, CK => CLK, Q => 
                           n21599, QN => n19234);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n4863, CK => CLK, Q => 
                           n21600, QN => n19235);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n4862, CK => CLK, Q => 
                           n21601, QN => n19236);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n4861, CK => CLK, Q => 
                           n21602, QN => n19237);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n4860, CK => CLK, Q => 
                           n21603, QN => n19238);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n4859, CK => CLK, Q => 
                           n21638, QN => n19239);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n4858, CK => CLK, Q => 
                           n21582, QN => n19240);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n4857, CK => CLK, Q => 
                           n21583, QN => n19241);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n4856, CK => CLK, Q => 
                           n21618, QN => n19242);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n4855, CK => CLK, Q => 
                           n21607, QN => n19243);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n4854, CK => CLK, Q => 
                           n21760, QN => n19244);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n4853, CK => CLK, Q => 
                           n21619, QN => n19245);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n4852, CK => CLK, Q => 
                           n21761, QN => n19246);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n4851, CK => CLK, Q => 
                           n21609, QN => n19247);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n4850, CK => CLK, Q => 
                           n21759, QN => n19248);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n4849, CK => CLK, Q => 
                           n21587, QN => n19249);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n4848, CK => CLK, Q => 
                           n21588, QN => n19250);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n4847, CK => CLK, Q => 
                           n21623, QN => n19251);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n4846, CK => CLK, Q => 
                           n21624, QN => n19252);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n4845, CK => CLK, Q => 
                           n21590, QN => n19253);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n4844, CK => CLK, Q => 
                           n21626, QN => n19254);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n4843, CK => CLK, Q => 
                           n21627, QN => n19255);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n4842, CK => CLK, Q => 
                           n21592, QN => n19256);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n4841, CK => CLK, Q => 
                           n21630, QN => n19257);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n4840, CK => CLK, Q => 
                           n21633, QN => n19258);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n4839, CK => CLK, Q => 
                           n21632, QN => n19259);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n4838, CK => CLK, Q => 
                           n21578, QN => n19260);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n4837, CK => CLK, Q => 
                           n21577, QN => n19261);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n4836, CK => CLK, Q => 
                           n21537, QN => n19262);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n4835, CK => CLK, Q => 
                           n21573, QN => n19263);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n4834, CK => CLK, Q => 
                           n21572, QN => n19264);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n4833, CK => CLK, Q => 
                           n21535, QN => n19265);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n4832, CK => CLK, Q => 
                           n21569, QN => n19266);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n4831, CK => CLK, Q => 
                           n21554, QN => n19267);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n4830, CK => CLK, Q => 
                           n21533, QN => n19268);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n4829, CK => CLK, Q => 
                           n21566, QN => n19269);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n4828, CK => CLK, Q => 
                           n21565, QN => n19270);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n4827, CK => CLK, Q => 
                           n21564, QN => n19271);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n4826, CK => CLK, Q => 
                           n21530, QN => n19272);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n4825, CK => CLK, Q => 
                           n21757, QN => n19273);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n4824, CK => CLK, Q => 
                           n21529, QN => n19274);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n4823, CK => CLK, Q => 
                           n21528, QN => n19275);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n4822, CK => CLK, Q => 
                           n21552, QN => n19276);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n4821, CK => CLK, Q => 
                           n21550, QN => n19277);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n4820, CK => CLK, Q => 
                           n21549, QN => n19278);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n4819, CK => CLK, Q => 
                           n21561, QN => n19279);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n4818, CK => CLK, Q => 
                           n21548, QN => n19280);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n4817, CK => CLK, Q => 
                           n21560, QN => n19281);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n4816, CK => CLK, Q => 
                           n21525, QN => n19282);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n4815, CK => CLK, Q => 
                           n21559, QN => n19283);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n4814, CK => CLK, Q => 
                           n21752, QN => n19284);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n4813, CK => CLK, Q => 
                           n21558, QN => n19285);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n4812, CK => CLK, Q => 
                           n21542, QN => n19286);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n4811, CK => CLK, Q => n21631
                           , QN => n19287);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n4810, CK => CLK, Q => n21555
                           , QN => n19288);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n4809, CK => CLK, Q => n21524
                           , QN => n19289);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n4808, CK => CLK, Q => n21539
                           , QN => n19290);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n4807, CK => CLK, Q => n21523
                           , QN => n19291);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n4806, CK => CLK, Q => n21841
                           , QN => n19292);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n4805, CK => CLK, Q => n21538
                           , QN => n19293);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n4804, CK => CLK, Q => n21540
                           , QN => n19294);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n4803, CK => CLK, Q => n21541
                           , QN => n19295);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n4802, CK => CLK, Q => n21556
                           , QN => n19296);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n4801, CK => CLK, Q => 
                           n21557, QN => n19297);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n4800, CK => CLK, Q => 
                           n21543, QN => n19298);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n4799, CK => CLK, Q => 
                           n21544, QN => n19299);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n4798, CK => CLK, Q => 
                           n21545, QN => n19300);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n4797, CK => CLK, Q => 
                           n21546, QN => n19301);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n4796, CK => CLK, Q => 
                           n21547, QN => n19302);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n4795, CK => CLK, Q => 
                           n21637, QN => n19303);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n4794, CK => CLK, Q => 
                           n21526, QN => n19304);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n4793, CK => CLK, Q => 
                           n21527, QN => n19305);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n4792, CK => CLK, Q => 
                           n21562, QN => n19306);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n4791, CK => CLK, Q => 
                           n21551, QN => n19307);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n4790, CK => CLK, Q => 
                           n21755, QN => n19308);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n4789, CK => CLK, Q => 
                           n21563, QN => n19309);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n4788, CK => CLK, Q => 
                           n21756, QN => n19310);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n4787, CK => CLK, Q => 
                           n21553, QN => n19311);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n4786, CK => CLK, Q => 
                           n21753, QN => n19312);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n4785, CK => CLK, Q => 
                           n21531, QN => n19313);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n4784, CK => CLK, Q => 
                           n21532, QN => n19314);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n4783, CK => CLK, Q => 
                           n21567, QN => n19315);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n4782, CK => CLK, Q => 
                           n21568, QN => n19316);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n4781, CK => CLK, Q => 
                           n21534, QN => n19317);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n4780, CK => CLK, Q => 
                           n21570, QN => n19318);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n4779, CK => CLK, Q => 
                           n21571, QN => n19319);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n4778, CK => CLK, Q => 
                           n21536, QN => n19320);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n4777, CK => CLK, Q => 
                           n21574, QN => n19321);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n4776, CK => CLK, Q => 
                           n21576, QN => n19322);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n4775, CK => CLK, Q => 
                           n21575, QN => n19323);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n4774, CK => CLK, Q => 
                           n21206, QN => n_1094);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n4773, CK => CLK, Q => 
                           n21205, QN => n_1095);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n4772, CK => CLK, Q => 
                           n21181, QN => n_1096);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n4771, CK => CLK, Q => 
                           n21173, QN => n_1097);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n4770, CK => CLK, Q => 
                           n21201, QN => n_1098);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n4769, CK => CLK, Q => 
                           n21179, QN => n_1099);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n4768, CK => CLK, Q => 
                           n21198, QN => n_1100);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n4767, CK => CLK, Q => 
                           n21192, QN => n_1101);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n4766, CK => CLK, Q => 
                           n21177, QN => n_1102);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n4765, CK => CLK, Q => 
                           n21197, QN => n_1103);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n4764, CK => CLK, Q => 
                           n21170, QN => n_1104);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n4763, CK => CLK, Q => 
                           n21169, QN => n_1105);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n4762, CK => CLK, Q => 
                           n21155, QN => n_1106);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n4761, CK => CLK, Q => 
                           n21277, QN => n_1107);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n4760, CK => CLK, Q => 
                           n21154, QN => n_1108);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n4759, CK => CLK, Q => 
                           n21153, QN => n_1109);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n4758, CK => CLK, Q => 
                           n21163, QN => n_1110);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n4757, CK => CLK, Q => 
                           n21189, QN => n_1111);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n4756, CK => CLK, Q => 
                           n21162, QN => n_1112);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n4755, CK => CLK, Q => 
                           n21195, QN => n_1113);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n4754, CK => CLK, Q => 
                           n21161, QN => n_1114);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n4753, CK => CLK, Q => 
                           n21167, QN => n_1115);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n4752, CK => CLK, Q => 
                           n21152, QN => n_1116);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n4751, CK => CLK, Q => 
                           n21166, QN => n_1117);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n4750, CK => CLK, Q => 
                           n21278, QN => n_1118);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n4749, CK => CLK, Q => 
                           n21194, QN => n_1119);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n4748, CK => CLK, Q => 
                           n21159, QN => n_1120);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n4747, CK => CLK, Q => 
                           n21207, QN => n_1121);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n4746, CK => CLK, Q => 
                           n21164, QN => n_1122);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n4745, CK => CLK, Q => 
                           n21174, QN => n_1123);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n4744, CK => CLK, Q => 
                           n21158, QN => n_1124);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n4743, CK => CLK, Q => 
                           n21151, QN => n_1125);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n4742, CK => CLK, Q => 
                           n21286, QN => n_1126);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n4741, CK => CLK, Q => 
                           n21182, QN => n_1127);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n4740, CK => CLK, Q => 
                           n21183, QN => n_1128);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n4739, CK => CLK, Q => 
                           n21184, QN => n_1129);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n4738, CK => CLK, Q => 
                           n21193, QN => n_1130);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n4737, CK => CLK, Q => 
                           n21165, QN => n_1131);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n4736, CK => CLK, Q => 
                           n21185, QN => n_1132);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n4735, CK => CLK, Q => 
                           n21186, QN => n_1133);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n4734, CK => CLK, Q => 
                           n21187, QN => n_1134);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n4733, CK => CLK, Q => 
                           n21160, QN => n_1135);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n4732, CK => CLK, Q => 
                           n21188, QN => n_1136);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n4731, CK => CLK, Q => 
                           n21209, QN => n_1137);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n4730, CK => CLK, Q => 
                           n21175, QN => n_1138);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n4729, CK => CLK, Q => 
                           n21176, QN => n_1139);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n4728, CK => CLK, Q => 
                           n21196, QN => n_1140);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n4727, CK => CLK, Q => 
                           n21190, QN => n_1141);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n4726, CK => CLK, Q => 
                           n21275, QN => n_1142);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n4725, CK => CLK, Q => 
                           n21168, QN => n_1143);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n4724, CK => CLK, Q => 
                           n21276, QN => n_1144);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n4723, CK => CLK, Q => 
                           n21191, QN => n_1145);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n4722, CK => CLK, Q => 
                           n21273, QN => n_1146);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n4721, CK => CLK, Q => 
                           n21156, QN => n_1147);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n4720, CK => CLK, Q => 
                           n21157, QN => n_1148);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n4719, CK => CLK, Q => 
                           n21171, QN => n_1149);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n4718, CK => CLK, Q => 
                           n21172, QN => n_1150);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n4717, CK => CLK, Q => 
                           n21178, QN => n_1151);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n4716, CK => CLK, Q => 
                           n21199, QN => n_1152);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n4715, CK => CLK, Q => 
                           n21200, QN => n_1153);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n4714, CK => CLK, Q => 
                           n21180, QN => n_1154);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n4713, CK => CLK, Q => 
                           n21202, QN => n_1155);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n4712, CK => CLK, Q => 
                           n21204, QN => n_1156);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n4711, CK => CLK, Q => 
                           n21203, QN => n_1157);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n4710, CK => CLK, Q => 
                           n21149, QN => n19388);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n4709, CK => CLK, Q => 
                           n21148, QN => n19389);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n4708, CK => CLK, Q => 
                           n21108, QN => n19390);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n4707, CK => CLK, Q => 
                           n21144, QN => n19391);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n4706, CK => CLK, Q => 
                           n21143, QN => n19392);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n4705, CK => CLK, Q => 
                           n21106, QN => n19393);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n4704, CK => CLK, Q => 
                           n21140, QN => n19394);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n4703, CK => CLK, Q => 
                           n21125, QN => n19395);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n4702, CK => CLK, Q => 
                           n21104, QN => n19396);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n4701, CK => CLK, Q => 
                           n21137, QN => n19397);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n4700, CK => CLK, Q => 
                           n21136, QN => n19398);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n4699, CK => CLK, Q => 
                           n21135, QN => n19399);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n4698, CK => CLK, Q => 
                           n21101, QN => n19400);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n4697, CK => CLK, Q => 
                           n21271, QN => n19401);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n4696, CK => CLK, Q => 
                           n21100, QN => n19402);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n4695, CK => CLK, Q => 
                           n21099, QN => n19403);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n4694, CK => CLK, Q => 
                           n21123, QN => n19404);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n4693, CK => CLK, Q => 
                           n21121, QN => n19405);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n4692, CK => CLK, Q => 
                           n21120, QN => n19406);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n4691, CK => CLK, Q => 
                           n21132, QN => n19407);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n4690, CK => CLK, Q => 
                           n21119, QN => n19408);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n4689, CK => CLK, Q => 
                           n21131, QN => n19409);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n4688, CK => CLK, Q => 
                           n21096, QN => n19410);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n4687, CK => CLK, Q => 
                           n21130, QN => n19411);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n4686, CK => CLK, Q => 
                           n21267, QN => n19412);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n4685, CK => CLK, Q => 
                           n21129, QN => n19413);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n4684, CK => CLK, Q => 
                           n21113, QN => n19414);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n4683, CK => CLK, Q => 
                           n21150, QN => n19415);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n4682, CK => CLK, Q => 
                           n21126, QN => n19416);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n4681, CK => CLK, Q => 
                           n21095, QN => n19417);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n4680, CK => CLK, Q => 
                           n21110, QN => n19418);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n4679, CK => CLK, Q => 
                           n21094, QN => n19419);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n4678, CK => CLK, Q => 
                           n21284, QN => n19420);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n4677, CK => CLK, Q => 
                           n21109, QN => n19421);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n4676, CK => CLK, Q => 
                           n21111, QN => n19422);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n4675, CK => CLK, Q => 
                           n21112, QN => n19423);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n4674, CK => CLK, Q => 
                           n21127, QN => n19424);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n4673, CK => CLK, Q => 
                           n21128, QN => n19425);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n4672, CK => CLK, Q => 
                           n21114, QN => n19426);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n4671, CK => CLK, Q => 
                           n21115, QN => n19427);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n4670, CK => CLK, Q => 
                           n21116, QN => n19428);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n4669, CK => CLK, Q => 
                           n21117, QN => n19429);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n4668, CK => CLK, Q => 
                           n21118, QN => n19430);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n4667, CK => CLK, Q => 
                           n21208, QN => n19431);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n4666, CK => CLK, Q => 
                           n21097, QN => n19432);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n4665, CK => CLK, Q => 
                           n21098, QN => n19433);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n4664, CK => CLK, Q => 
                           n21133, QN => n19434);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n4663, CK => CLK, Q => 
                           n21122, QN => n19435);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n4662, CK => CLK, Q => 
                           n21269, QN => n19436);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n4661, CK => CLK, Q => 
                           n21134, QN => n19437);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n4660, CK => CLK, Q => 
                           n21270, QN => n19438);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n4659, CK => CLK, Q => 
                           n21124, QN => n19439);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n4658, CK => CLK, Q => 
                           n21268, QN => n19440);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n4657, CK => CLK, Q => 
                           n21102, QN => n19441);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n4656, CK => CLK, Q => 
                           n21103, QN => n19442);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n4655, CK => CLK, Q => 
                           n21138, QN => n19443);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n4654, CK => CLK, Q => 
                           n21139, QN => n19444);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n4653, CK => CLK, Q => 
                           n21105, QN => n19445);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n4652, CK => CLK, Q => 
                           n21141, QN => n19446);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n4651, CK => CLK, Q => 
                           n21142, QN => n19447);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n4650, CK => CLK, Q => 
                           n21107, QN => n19448);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n4649, CK => CLK, Q => 
                           n21145, QN => n19449);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n4648, CK => CLK, Q => 
                           n21147, QN => n19450);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n4647, CK => CLK, Q => 
                           n21146, QN => n19451);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n4646, CK => CLK, Q => 
                           n22223, QN => n19452);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n4645, CK => CLK, Q => 
                           n22222, QN => n19453);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n4644, CK => CLK, Q => 
                           n22220, QN => n19454);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n4643, CK => CLK, Q => 
                           n22084, QN => n19455);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n4642, CK => CLK, Q => 
                           n22217, QN => n19456);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n4641, CK => CLK, Q => 
                           n22215, QN => n19457);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n4640, CK => CLK, Q => 
                           n22213, QN => n19458);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n4639, CK => CLK, Q => 
                           n22211, QN => n19459);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n4638, CK => CLK, Q => 
                           n22210, QN => n19460);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n4637, CK => CLK, Q => 
                           n22209, QN => n19461);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n4636, CK => CLK, Q => 
                           n22080, QN => n19462);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n4635, CK => CLK, Q => 
                           n22078, QN => n19463);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n4634, CK => CLK, Q => 
                           n22076, QN => n19464);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n4633, CK => CLK, Q => 
                           n22075, QN => n19465);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n4632, CK => CLK, Q => 
                           n22073, QN => n19466);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n4631, CK => CLK, Q => 
                           n22071, QN => n19467);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n4630, CK => CLK, Q => 
                           n22069, QN => n19468);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n4629, CK => CLK, Q => 
                           n22206, QN => n19469);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n4628, CK => CLK, Q => 
                           n22068, QN => n19470);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n4627, CK => CLK, Q => 
                           n22203, QN => n19471);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n4626, CK => CLK, Q => 
                           n22067, QN => n19472);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n4625, CK => CLK, Q => 
                           n22066, QN => n19473);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n4624, CK => CLK, Q => 
                           n22065, QN => n19474);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n4623, CK => CLK, Q => 
                           n22063, QN => n19475);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n4622, CK => CLK, Q => 
                           n22199, QN => n19476);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n4621, CK => CLK, Q => 
                           n22197, QN => n19477);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n4620, CK => CLK, Q => 
                           n22062, QN => n19478);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n4619, CK => CLK, Q => 
                           n22195, QN => n19479);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n4618, CK => CLK, Q => 
                           n22060, QN => n19480);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n4617, CK => CLK, Q => 
                           n22192, QN => n19481);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n4616, CK => CLK, Q => 
                           n22059, QN => n19482);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n4615, CK => CLK, Q => 
                           n22058, QN => n19483);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n4614, CK => CLK, Q => 
                           n22225, QN => n19484);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n4613, CK => CLK, Q => 
                           n22190, QN => n19485);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n4612, CK => CLK, Q => 
                           n22191, QN => n19486);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n4611, CK => CLK, Q => 
                           n22193, QN => n19487);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n4610, CK => CLK, Q => 
                           n22194, QN => n19488);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n4609, CK => CLK, Q => 
                           n22061, QN => n19489);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n4608, CK => CLK, Q => 
                           n22196, QN => n19490);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n4607, CK => CLK, Q => 
                           n22198, QN => n19491);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n4606, CK => CLK, Q => 
                           n22200, QN => n19492);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n4605, CK => CLK, Q => 
                           n22064, QN => n19493);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n4604, CK => CLK, Q => 
                           n22201, QN => n19494);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n4603, CK => CLK, Q => 
                           n22086, QN => n19495);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n4602, CK => CLK, Q => 
                           n22202, QN => n19496);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n4601, CK => CLK, Q => 
                           n22204, QN => n19497);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n4600, CK => CLK, Q => 
                           n22205, QN => n19498);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n4599, CK => CLK, Q => 
                           n22207, QN => n19499);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n4598, CK => CLK, Q => 
                           n22070, QN => n19500);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n4597, CK => CLK, Q => 
                           n22072, QN => n19501);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n4596, CK => CLK, Q => 
                           n22074, QN => n19502);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n4595, CK => CLK, Q => 
                           n22208, QN => n19503);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n4594, CK => CLK, Q => 
                           n22077, QN => n19504);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n4593, CK => CLK, Q => 
                           n22079, QN => n19505);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n4592, CK => CLK, Q => 
                           n22081, QN => n19506);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n4591, CK => CLK, Q => 
                           n22082, QN => n19507);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n4590, CK => CLK, Q => 
                           n22083, QN => n19508);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n4589, CK => CLK, Q => 
                           n22212, QN => n19509);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n4588, CK => CLK, Q => 
                           n22214, QN => n19510);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n4587, CK => CLK, Q => 
                           n22216, QN => n19511);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n4586, CK => CLK, Q => 
                           n22218, QN => n19512);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n4585, CK => CLK, Q => 
                           n22219, QN => n19513);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n4584, CK => CLK, Q => 
                           n22221, QN => n19514);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n4583, CK => CLK, Q => 
                           n22085, QN => n19515);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n4582, CK => CLK, Q => 
                           n22336, QN => n19516);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n4581, CK => CLK, Q => 
                           n22397, QN => n19517);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n4580, CK => CLK, Q => 
                           n22337, QN => n19518);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n4579, CK => CLK, Q => 
                           n22358, QN => n19519);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n4578, CK => CLK, Q => 
                           n22338, QN => n19520);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n4577, CK => CLK, Q => 
                           n22292, QN => n19521);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n4576, CK => CLK, Q => 
                           n22293, QN => n19522);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n4575, CK => CLK, Q => 
                           n22294, QN => n19523);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n4574, CK => CLK, Q => 
                           n22295, QN => n19524);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n4573, CK => CLK, Q => 
                           n22296, QN => n19525);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n4572, CK => CLK, Q => 
                           n22339, QN => n19526);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n4571, CK => CLK, Q => 
                           n22340, QN => n19527);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n4570, CK => CLK, Q => 
                           n22341, QN => n19528);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n4569, CK => CLK, Q => 
                           n22342, QN => n19529);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n4568, CK => CLK, Q => 
                           n22380, QN => n19530);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n4567, CK => CLK, Q => 
                           n22359, QN => n19531);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n4566, CK => CLK, Q => 
                           n22343, QN => n19532);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n4565, CK => CLK, Q => 
                           n22297, QN => n19533);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n4564, CK => CLK, Q => 
                           n22298, QN => n19534);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n4563, CK => CLK, Q => 
                           n22299, QN => n19535);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n4562, CK => CLK, Q => 
                           n22300, QN => n19536);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n4561, CK => CLK, Q => 
                           n22344, QN => n19537);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n4560, CK => CLK, Q => 
                           n22398, QN => n19538);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n4559, CK => CLK, Q => 
                           n22399, QN => n19539);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n4558, CK => CLK, Q => 
                           n22348, QN => n19540);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n4557, CK => CLK, Q => 
                           n22349, QN => n19541);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n4556, CK => CLK, Q => 
                           n22350, QN => n19542);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n4555, CK => CLK, Q => 
                           n22351, QN => n19543);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n4554, CK => CLK, Q => 
                           n22301, QN => n19544);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n4553, CK => CLK, Q => 
                           n22352, QN => n19545);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n4552, CK => CLK, Q => 
                           n22345, QN => n19546);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n4551, CK => CLK, Q => 
                           n22302, QN => n19547);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n4550, CK => CLK, Q => 
                           n22290, QN => n19548);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n4549, CK => CLK, Q => 
                           n22303, QN => n19549);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n4548, CK => CLK, Q => 
                           n22304, QN => n19550);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n4547, CK => CLK, Q => 
                           n22353, QN => n19551);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n4546, CK => CLK, Q => 
                           n22354, QN => n19552);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n4545, CK => CLK, Q => 
                           n22360, QN => n19553);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n4544, CK => CLK, Q => 
                           n22355, QN => n19554);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n4543, CK => CLK, Q => 
                           n22356, QN => n19555);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n4542, CK => CLK, Q => 
                           n22357, QN => n19556);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n4541, CK => CLK, Q => 
                           n22305, QN => n19557);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n4540, CK => CLK, Q => 
                           n22306, QN => n19558);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n4539, CK => CLK, Q => 
                           n22482, QN => n19559);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n4538, CK => CLK, Q => 
                           n22346, QN => n19560);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n4537, CK => CLK, Q => 
                           n22361, QN => n19561);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n4536, CK => CLK, Q => 
                           n22362, QN => n19562);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n4535, CK => CLK, Q => 
                           n22400, QN => n19563);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n4534, CK => CLK, Q => 
                           n22363, QN => n19564);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n4533, CK => CLK, Q => 
                           n22364, QN => n19565);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n4532, CK => CLK, Q => 
                           n22381, QN => n19566);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n4531, CK => CLK, Q => 
                           n22365, QN => n19567);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n4530, CK => CLK, Q => 
                           n22347, QN => n19568);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n4529, CK => CLK, Q => 
                           n22307, QN => n19569);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n4528, CK => CLK, Q => 
                           n22308, QN => n19570);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n4527, CK => CLK, Q => 
                           n22309, QN => n19571);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n4526, CK => CLK, Q => 
                           n22310, QN => n19572);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n4525, CK => CLK, Q => 
                           n22366, QN => n19573);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n4524, CK => CLK, Q => 
                           n22368, QN => n19574);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n4523, CK => CLK, Q => 
                           n22369, QN => n19575);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n4522, CK => CLK, Q => 
                           n22401, QN => n19576);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n4521, CK => CLK, Q => 
                           n22370, QN => n19577);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n4520, CK => CLK, Q => 
                           n22410, QN => n19578);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n4519, CK => CLK, Q => 
                           n22371, QN => n19579);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n4518, CK => CLK, Q => 
                           n22142, QN => n19580);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n4517, CK => CLK, Q => 
                           n22140, QN => n19581);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n4516, CK => CLK, Q => 
                           n22138, QN => n19582);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n4515, CK => CLK, Q => 
                           n22136, QN => n19583);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n4514, CK => CLK, Q => 
                           n22134, QN => n19584);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n4513, CK => CLK, Q => 
                           n22132, QN => n19585);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n4512, CK => CLK, Q => 
                           n22130, QN => n19586);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n4511, CK => CLK, Q => 
                           n22128, QN => n19587);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n4510, CK => CLK, Q => 
                           n22126, QN => n19588);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n4509, CK => CLK, Q => 
                           n22124, QN => n19589);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n4508, CK => CLK, Q => 
                           n22122, QN => n19590);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n4507, CK => CLK, Q => 
                           n22120, QN => n19591);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n4506, CK => CLK, Q => 
                           n22119, QN => n19592);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n4505, CK => CLK, Q => 
                           n22188, QN => n19593);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n4504, CK => CLK, Q => 
                           n22117, QN => n19594);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n4503, CK => CLK, Q => 
                           n22115, QN => n19595);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n4502, CK => CLK, Q => 
                           n22114, QN => n19596);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n4501, CK => CLK, Q => 
                           n22112, QN => n19597);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n4500, CK => CLK, Q => 
                           n22110, QN => n19598);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n4499, CK => CLK, Q => 
                           n22108, QN => n19599);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n4498, CK => CLK, Q => 
                           n22106, QN => n19600);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n4497, CK => CLK, Q => 
                           n22105, QN => n19601);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n4496, CK => CLK, Q => 
                           n22103, QN => n19602);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n4495, CK => CLK, Q => 
                           n22101, QN => n19603);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n4494, CK => CLK, Q => 
                           n22185, QN => n19604);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n4493, CK => CLK, Q => 
                           n22098, QN => n19605);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n4492, CK => CLK, Q => 
                           n22096, QN => n19606);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n4491, CK => CLK, Q => 
                           n22184, QN => n19607);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n4490, CK => CLK, Q => 
                           n22093, QN => n19608);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n4489, CK => CLK, Q => 
                           n22091, QN => n19609);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n4488, CK => CLK, Q => 
                           n22089, QN => n19610);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n4487, CK => CLK, Q => 
                           n22087, QN => n19611);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n4486, CK => CLK, Q => 
                           n22417, QN => n19612);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n4485, CK => CLK, Q => 
                           n22088, QN => n19613);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n4484, CK => CLK, Q => 
                           n22090, QN => n19614);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n4483, CK => CLK, Q => 
                           n22092, QN => n19615);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n4482, CK => CLK, Q => 
                           n22094, QN => n19616);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n4481, CK => CLK, Q => 
                           n22095, QN => n19617);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n4480, CK => CLK, Q => 
                           n22097, QN => n19618);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n4479, CK => CLK, Q => 
                           n22099, QN => n19619);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n4478, CK => CLK, Q => 
                           n22100, QN => n19620);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n4477, CK => CLK, Q => 
                           n22102, QN => n19621);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n4476, CK => CLK, Q => 
                           n22104, QN => n19622);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n4475, CK => CLK, Q => 
                           n22224, QN => n19623);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n4474, CK => CLK, Q => 
                           n22107, QN => n19624);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n4473, CK => CLK, Q => 
                           n22109, QN => n19625);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n4472, CK => CLK, Q => 
                           n22111, QN => n19626);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n4471, CK => CLK, Q => 
                           n22113, QN => n19627);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n4470, CK => CLK, Q => 
                           n22186, QN => n19628);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n4469, CK => CLK, Q => 
                           n22116, QN => n19629);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n4468, CK => CLK, Q => 
                           n22187, QN => n19630);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n4467, CK => CLK, Q => 
                           n22118, QN => n19631);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n4466, CK => CLK, Q => 
                           n22189, QN => n19632);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n4465, CK => CLK, Q => 
                           n22121, QN => n19633);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n4464, CK => CLK, Q => 
                           n22123, QN => n19634);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n4463, CK => CLK, Q => 
                           n22125, QN => n19635);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n4462, CK => CLK, Q => 
                           n22127, QN => n19636);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n4461, CK => CLK, Q => 
                           n22129, QN => n19637);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n4460, CK => CLK, Q => 
                           n22131, QN => n19638);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n4459, CK => CLK, Q => 
                           n22133, QN => n19639);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n4458, CK => CLK, Q => 
                           n22135, QN => n19640);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n4457, CK => CLK, Q => 
                           n22137, QN => n19641);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n4456, CK => CLK, Q => 
                           n22139, QN => n19642);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n4455, CK => CLK, Q => 
                           n22141, QN => n19643);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n4454, CK => CLK, Q => 
                           n22373, QN => n19644);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n4453, CK => CLK, Q => 
                           n22374, QN => n19645);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n4452, CK => CLK, Q => 
                           n22375, QN => n19646);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n4451, CK => CLK, Q => 
                           n22376, QN => n19647);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n4450, CK => CLK, Q => 
                           n22367, QN => n19648);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n4449, CK => CLK, Q => 
                           n22311, QN => n19649);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n4448, CK => CLK, Q => 
                           n22312, QN => n19650);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n4447, CK => CLK, Q => 
                           n22313, QN => n19651);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n4446, CK => CLK, Q => 
                           n22314, QN => n19652);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n4445, CK => CLK, Q => 
                           n22315, QN => n19653);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n4444, CK => CLK, Q => 
                           n22377, QN => n19654);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n4443, CK => CLK, Q => 
                           n22382, QN => n19655);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n4442, CK => CLK, Q => 
                           n22383, QN => n19656);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n4441, CK => CLK, Q => 
                           n22384, QN => n19657);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n4440, CK => CLK, Q => 
                           n22385, QN => n19658);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n4439, CK => CLK, Q => 
                           n22386, QN => n19659);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n4438, CK => CLK, Q => 
                           n22316, QN => n19660);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n4437, CK => CLK, Q => 
                           n22317, QN => n19661);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n4436, CK => CLK, Q => 
                           n22318, QN => n19662);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n4435, CK => CLK, Q => 
                           n22319, QN => n19663);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n4434, CK => CLK, Q => 
                           n22320, QN => n19664);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n4433, CK => CLK, Q => 
                           n22378, QN => n19665);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n4432, CK => CLK, Q => 
                           n22321, QN => n19666);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n4431, CK => CLK, Q => 
                           n22387, QN => n19667);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n4430, CK => CLK, Q => 
                           n22388, QN => n19668);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n4429, CK => CLK, Q => 
                           n22402, QN => n19669);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n4428, CK => CLK, Q => 
                           n22389, QN => n19670);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n4427, CK => CLK, Q => 
                           n22390, QN => n19671);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n4426, CK => CLK, Q => 
                           n22322, QN => n19672);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n4425, CK => CLK, Q => 
                           n22323, QN => n19673);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n4424, CK => CLK, Q => 
                           n22324, QN => n19674);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n4423, CK => CLK, Q => 
                           n22325, QN => n19675);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n4422, CK => CLK, Q => 
                           n22372, QN => n19676);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n4421, CK => CLK, Q => 
                           n22326, QN => n19677);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n4420, CK => CLK, Q => 
                           n22379, QN => n19678);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n4419, CK => CLK, Q => 
                           n22391, QN => n19679);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n4418, CK => CLK, Q => 
                           n22392, QN => n19680);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n4417, CK => CLK, Q => 
                           n22393, QN => n19681);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n4416, CK => CLK, Q => 
                           n22394, QN => n19682);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n4415, CK => CLK, Q => 
                           n22395, QN => n19683);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n4414, CK => CLK, Q => 
                           n22327, QN => n19684);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n4413, CK => CLK, Q => 
                           n22328, QN => n19685);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n4412, CK => CLK, Q => 
                           n22329, QN => n19686);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n4411, CK => CLK, Q => 
                           n22483, QN => n19687);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n4410, CK => CLK, Q => 
                           n22330, QN => n19688);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n4409, CK => CLK, Q => 
                           n22396, QN => n19689);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n4408, CK => CLK, Q => 
                           n22403, QN => n19690);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n4407, CK => CLK, Q => 
                           n22404, QN => n19691);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n4406, CK => CLK, Q => 
                           n22405, QN => n19692);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n4405, CK => CLK, Q => 
                           n22406, QN => n19693);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n4404, CK => CLK, Q => 
                           n22407, QN => n19694);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n4403, CK => CLK, Q => 
                           n22408, QN => n19695);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n4402, CK => CLK, Q => 
                           n22331, QN => n19696);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n4401, CK => CLK, Q => 
                           n22332, QN => n19697);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n4400, CK => CLK, Q => 
                           n22333, QN => n19698);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n4399, CK => CLK, Q => 
                           n22334, QN => n19699);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n4398, CK => CLK, Q => 
                           n22335, QN => n19700);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n4397, CK => CLK, Q => 
                           n22409, QN => n19701);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n4396, CK => CLK, Q => 
                           n22411, QN => n19702);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n4395, CK => CLK, Q => 
                           n22412, QN => n19703);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n4394, CK => CLK, Q => 
                           n22413, QN => n19704);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n4393, CK => CLK, Q => 
                           n22414, QN => n19705);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n4392, CK => CLK, Q => 
                           n22415, QN => n19706);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n4391, CK => CLK, Q => 
                           n22416, QN => n19707);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n4390, CK => CLK, Q => 
                           n_1158, QN => n19708);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n4389, CK => CLK, Q => 
                           n_1159, QN => n19709);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n4388, CK => CLK, Q => 
                           n_1160, QN => n19710);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n4387, CK => CLK, Q => 
                           n_1161, QN => n19711);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n4386, CK => CLK, Q => 
                           n_1162, QN => n19712);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n4385, CK => CLK, Q => 
                           n_1163, QN => n19713);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n4384, CK => CLK, Q => 
                           n_1164, QN => n19714);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n4383, CK => CLK, Q => 
                           n_1165, QN => n19715);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n4382, CK => CLK, Q => 
                           n_1166, QN => n19716);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n4381, CK => CLK, Q => 
                           n_1167, QN => n19717);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n4380, CK => CLK, Q => 
                           n_1168, QN => n19718);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n4379, CK => CLK, Q => 
                           n_1169, QN => n19719);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n4378, CK => CLK, Q => 
                           n_1170, QN => n19720);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n4377, CK => CLK, Q => 
                           n_1171, QN => n19721);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n4376, CK => CLK, Q => 
                           n_1172, QN => n19722);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n4375, CK => CLK, Q => 
                           n_1173, QN => n19723);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n4374, CK => CLK, Q => 
                           n_1174, QN => n19724);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n4373, CK => CLK, Q => 
                           n_1175, QN => n19725);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n4372, CK => CLK, Q => 
                           n_1176, QN => n19726);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n4371, CK => CLK, Q => 
                           n_1177, QN => n19727);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n4370, CK => CLK, Q => 
                           n_1178, QN => n19728);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n4369, CK => CLK, Q => 
                           n_1179, QN => n19729);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n4368, CK => CLK, Q => 
                           n_1180, QN => n19730);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n4367, CK => CLK, Q => 
                           n_1181, QN => n19731);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n4366, CK => CLK, Q => 
                           n_1182, QN => n19732);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n4365, CK => CLK, Q => 
                           n_1183, QN => n19733);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n4364, CK => CLK, Q => 
                           n_1184, QN => n19734);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n4363, CK => CLK, Q => 
                           n_1185, QN => n19735);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n4362, CK => CLK, Q => 
                           n_1186, QN => n19736);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n4361, CK => CLK, Q => 
                           n_1187, QN => n19737);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n4360, CK => CLK, Q => 
                           n_1188, QN => n19738);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n4359, CK => CLK, Q => 
                           n_1189, QN => n19739);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n4358, CK => CLK, Q => 
                           n_1190, QN => n19740);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n4357, CK => CLK, Q => 
                           n_1191, QN => n19741);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n4356, CK => CLK, Q => 
                           n_1192, QN => n19742);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n4355, CK => CLK, Q => 
                           n_1193, QN => n19743);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n4354, CK => CLK, Q => 
                           n_1194, QN => n19744);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n4353, CK => CLK, Q => 
                           n_1195, QN => n19745);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n4352, CK => CLK, Q => 
                           n_1196, QN => n19746);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n4351, CK => CLK, Q => 
                           n_1197, QN => n19747);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n4350, CK => CLK, Q => 
                           n_1198, QN => n19748);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n4349, CK => CLK, Q => 
                           n_1199, QN => n19749);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n4348, CK => CLK, Q => 
                           n_1200, QN => n19750);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n4347, CK => CLK, Q => 
                           n_1201, QN => n19751);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n4346, CK => CLK, Q => 
                           n_1202, QN => n19752);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n4345, CK => CLK, Q => 
                           n_1203, QN => n19753);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n4344, CK => CLK, Q => 
                           n_1204, QN => n19754);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n4343, CK => CLK, Q => 
                           n_1205, QN => n19755);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n4342, CK => CLK, Q => 
                           n_1206, QN => n19756);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n4341, CK => CLK, Q => 
                           n_1207, QN => n19757);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n4340, CK => CLK, Q => 
                           n_1208, QN => n19758);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n4339, CK => CLK, Q => 
                           n_1209, QN => n19759);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n4338, CK => CLK, Q => 
                           n_1210, QN => n19760);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n4337, CK => CLK, Q => 
                           n_1211, QN => n19761);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n4336, CK => CLK, Q => 
                           n_1212, QN => n19762);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n4335, CK => CLK, Q => 
                           n_1213, QN => n19763);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n4334, CK => CLK, Q => 
                           n_1214, QN => n19764);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n4333, CK => CLK, Q => 
                           n_1215, QN => n19765);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n4332, CK => CLK, Q => 
                           n_1216, QN => n19766);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n4331, CK => CLK, Q => 
                           n_1217, QN => n19767);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n4330, CK => CLK, Q => 
                           n_1218, QN => n19768);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n4329, CK => CLK, Q => 
                           n_1219, QN => n19769);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n4328, CK => CLK, Q => 
                           n_1220, QN => n19770);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n4327, CK => CLK, Q => 
                           n_1221, QN => n19771);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n4326, CK => CLK, Q => 
                           n_1222, QN => n19772);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n4325, CK => CLK, Q => 
                           n_1223, QN => n19773);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n4324, CK => CLK, Q => 
                           n_1224, QN => n19774);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n4323, CK => CLK, Q => 
                           n_1225, QN => n19775);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n4322, CK => CLK, Q => 
                           n_1226, QN => n19776);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n4321, CK => CLK, Q => 
                           n_1227, QN => n19777);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n4320, CK => CLK, Q => 
                           n_1228, QN => n19778);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n4319, CK => CLK, Q => 
                           n_1229, QN => n19779);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n4318, CK => CLK, Q => 
                           n_1230, QN => n19780);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n4317, CK => CLK, Q => 
                           n_1231, QN => n19781);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n4316, CK => CLK, Q => 
                           n_1232, QN => n19782);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n4315, CK => CLK, Q => 
                           n_1233, QN => n19783);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n4314, CK => CLK, Q => 
                           n_1234, QN => n19784);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n4313, CK => CLK, Q => 
                           n_1235, QN => n19785);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n4312, CK => CLK, Q => 
                           n_1236, QN => n19786);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n4311, CK => CLK, Q => 
                           n_1237, QN => n19787);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n4310, CK => CLK, Q => 
                           n_1238, QN => n19788);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n4309, CK => CLK, Q => 
                           n_1239, QN => n19789);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n4308, CK => CLK, Q => 
                           n_1240, QN => n19790);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n4307, CK => CLK, Q => 
                           n_1241, QN => n19791);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n4306, CK => CLK, Q => 
                           n_1242, QN => n19792);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n4305, CK => CLK, Q => 
                           n_1243, QN => n19793);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n4304, CK => CLK, Q => 
                           n_1244, QN => n19794);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n4303, CK => CLK, Q => 
                           n_1245, QN => n19795);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n4302, CK => CLK, Q => 
                           n_1246, QN => n19796);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n4301, CK => CLK, Q => 
                           n_1247, QN => n19797);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n4300, CK => CLK, Q => 
                           n_1248, QN => n19798);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n4299, CK => CLK, Q => 
                           n_1249, QN => n19799);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n4298, CK => CLK, Q => 
                           n_1250, QN => n19800);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n4297, CK => CLK, Q => 
                           n_1251, QN => n19801);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n4296, CK => CLK, Q => 
                           n_1252, QN => n19802);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n4295, CK => CLK, Q => 
                           n_1253, QN => n19803);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n4294, CK => CLK, Q => 
                           n_1254, QN => n19804);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n4293, CK => CLK, Q => 
                           n_1255, QN => n19805);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n4292, CK => CLK, Q => 
                           n_1256, QN => n19806);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n4291, CK => CLK, Q => 
                           n_1257, QN => n19807);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n4290, CK => CLK, Q => 
                           n_1258, QN => n19808);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n4289, CK => CLK, Q => 
                           n_1259, QN => n19809);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n4288, CK => CLK, Q => 
                           n_1260, QN => n19810);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n4287, CK => CLK, Q => 
                           n_1261, QN => n19811);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n4286, CK => CLK, Q => 
                           n_1262, QN => n19812);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n4285, CK => CLK, Q => 
                           n_1263, QN => n19813);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n4284, CK => CLK, Q => 
                           n_1264, QN => n19814);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n4283, CK => CLK, Q => 
                           n_1265, QN => n19815);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n4282, CK => CLK, Q => 
                           n_1266, QN => n19816);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n4281, CK => CLK, Q => 
                           n_1267, QN => n19817);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n4280, CK => CLK, Q => 
                           n_1268, QN => n19818);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n4279, CK => CLK, Q => 
                           n_1269, QN => n19819);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n4278, CK => CLK, Q => 
                           n_1270, QN => n19820);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n4277, CK => CLK, Q => 
                           n_1271, QN => n19821);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n4276, CK => CLK, Q => 
                           n_1272, QN => n19822);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n4275, CK => CLK, Q => 
                           n_1273, QN => n19823);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n4274, CK => CLK, Q => 
                           n_1274, QN => n19824);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n4273, CK => CLK, Q => 
                           n_1275, QN => n19825);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n4272, CK => CLK, Q => 
                           n_1276, QN => n19826);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n4271, CK => CLK, Q => 
                           n_1277, QN => n19827);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n4270, CK => CLK, Q => 
                           n_1278, QN => n19828);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n4269, CK => CLK, Q => 
                           n_1279, QN => n19829);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n4268, CK => CLK, Q => 
                           n_1280, QN => n19830);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n4267, CK => CLK, Q => 
                           n_1281, QN => n19831);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n4266, CK => CLK, Q => 
                           n_1282, QN => n19832);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n4265, CK => CLK, Q => 
                           n_1283, QN => n19833);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n4264, CK => CLK, Q => 
                           n_1284, QN => n19834);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n4263, CK => CLK, Q => 
                           n_1285, QN => n19835);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n4262, CK => CLK, Q => 
                           n_1286, QN => n19836);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n4261, CK => CLK, Q => 
                           n_1287, QN => n19837);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n4260, CK => CLK, Q => 
                           n_1288, QN => n19838);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n4259, CK => CLK, Q => 
                           n_1289, QN => n19839);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n4258, CK => CLK, Q => 
                           n_1290, QN => n19840);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n4257, CK => CLK, Q => 
                           n_1291, QN => n19841);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n4256, CK => CLK, Q => 
                           n_1292, QN => n19842);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n4255, CK => CLK, Q => 
                           n_1293, QN => n19843);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n4254, CK => CLK, Q => 
                           n_1294, QN => n19844);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n4253, CK => CLK, Q => 
                           n_1295, QN => n19845);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n4252, CK => CLK, Q => 
                           n_1296, QN => n19846);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n4251, CK => CLK, Q => 
                           n_1297, QN => n19847);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n4250, CK => CLK, Q => 
                           n_1298, QN => n19848);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n4249, CK => CLK, Q => 
                           n_1299, QN => n19849);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n4248, CK => CLK, Q => 
                           n_1300, QN => n19850);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n4247, CK => CLK, Q => 
                           n_1301, QN => n19851);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n4246, CK => CLK, Q => 
                           n_1302, QN => n19852);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n4245, CK => CLK, Q => 
                           n_1303, QN => n19853);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n4244, CK => CLK, Q => 
                           n_1304, QN => n19854);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n4243, CK => CLK, Q => 
                           n_1305, QN => n19855);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n4242, CK => CLK, Q => 
                           n_1306, QN => n19856);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n4241, CK => CLK, Q => 
                           n_1307, QN => n19857);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n4240, CK => CLK, Q => 
                           n_1308, QN => n19858);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n4239, CK => CLK, Q => 
                           n_1309, QN => n19859);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n4238, CK => CLK, Q => 
                           n_1310, QN => n19860);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n4237, CK => CLK, Q => 
                           n_1311, QN => n19861);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n4236, CK => CLK, Q => 
                           n_1312, QN => n19862);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n4235, CK => CLK, Q => 
                           n_1313, QN => n19863);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n4234, CK => CLK, Q => 
                           n_1314, QN => n19864);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n4233, CK => CLK, Q => 
                           n_1315, QN => n19865);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n4232, CK => CLK, Q => 
                           n_1316, QN => n19866);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n4231, CK => CLK, Q => 
                           n_1317, QN => n19867);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n4230, CK => CLK, Q => 
                           n_1318, QN => n19868);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n4229, CK => CLK, Q => 
                           n_1319, QN => n19869);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n4228, CK => CLK, Q => 
                           n_1320, QN => n19870);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n4227, CK => CLK, Q => 
                           n_1321, QN => n19871);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n4226, CK => CLK, Q => 
                           n_1322, QN => n19872);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n4225, CK => CLK, Q => 
                           n_1323, QN => n19873);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n4224, CK => CLK, Q => 
                           n_1324, QN => n19874);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n4223, CK => CLK, Q => 
                           n_1325, QN => n19875);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n4222, CK => CLK, Q => 
                           n_1326, QN => n19876);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n4221, CK => CLK, Q => 
                           n_1327, QN => n19877);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n4220, CK => CLK, Q => 
                           n_1328, QN => n19878);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n4219, CK => CLK, Q => 
                           n_1329, QN => n19879);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n4218, CK => CLK, Q => 
                           n_1330, QN => n19880);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n4217, CK => CLK, Q => 
                           n_1331, QN => n19881);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n4216, CK => CLK, Q => 
                           n_1332, QN => n19882);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n4215, CK => CLK, Q => 
                           n_1333, QN => n19883);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n4214, CK => CLK, Q => 
                           n_1334, QN => n19884);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n4213, CK => CLK, Q => 
                           n_1335, QN => n19885);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n4212, CK => CLK, Q => 
                           n_1336, QN => n19886);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n4211, CK => CLK, Q => 
                           n_1337, QN => n19887);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n4210, CK => CLK, Q => 
                           n_1338, QN => n19888);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n4209, CK => CLK, Q => 
                           n_1339, QN => n19889);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n4208, CK => CLK, Q => 
                           n_1340, QN => n19890);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n4207, CK => CLK, Q => 
                           n_1341, QN => n19891);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n4206, CK => CLK, Q => 
                           n_1342, QN => n19892);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n4205, CK => CLK, Q => 
                           n_1343, QN => n19893);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n4204, CK => CLK, Q => 
                           n_1344, QN => n19894);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n4203, CK => CLK, Q => 
                           n_1345, QN => n19895);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n4202, CK => CLK, Q => 
                           n_1346, QN => n19896);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n4201, CK => CLK, Q => 
                           n_1347, QN => n19897);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n4200, CK => CLK, Q => 
                           n_1348, QN => n19898);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n4199, CK => CLK, Q => 
                           n_1349, QN => n19899);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n4198, CK => CLK, Q => 
                           n_1350, QN => n19900);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n4197, CK => CLK, Q => 
                           n_1351, QN => n19901);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n4196, CK => CLK, Q => 
                           n_1352, QN => n19902);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n4195, CK => CLK, Q => 
                           n_1353, QN => n19903);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n4194, CK => CLK, Q => 
                           n_1354, QN => n19904);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n4193, CK => CLK, Q => 
                           n_1355, QN => n19905);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n4192, CK => CLK, Q => 
                           n_1356, QN => n19906);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n4191, CK => CLK, Q => 
                           n_1357, QN => n19907);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n4190, CK => CLK, Q => 
                           n_1358, QN => n19908);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n4189, CK => CLK, Q => 
                           n_1359, QN => n19909);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n4188, CK => CLK, Q => 
                           n_1360, QN => n19910);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n4187, CK => CLK, Q => 
                           n_1361, QN => n19911);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n4186, CK => CLK, Q => 
                           n_1362, QN => n19912);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n4185, CK => CLK, Q => 
                           n_1363, QN => n19913);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n4184, CK => CLK, Q => 
                           n_1364, QN => n19914);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n4183, CK => CLK, Q => 
                           n_1365, QN => n19915);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n4182, CK => CLK, Q => 
                           n_1366, QN => n19916);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n4181, CK => CLK, Q => 
                           n_1367, QN => n19917);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n4180, CK => CLK, Q => 
                           n_1368, QN => n19918);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n4179, CK => CLK, Q => 
                           n_1369, QN => n19919);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n4178, CK => CLK, Q => 
                           n_1370, QN => n19920);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n4177, CK => CLK, Q => 
                           n_1371, QN => n19921);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n4176, CK => CLK, Q => 
                           n_1372, QN => n19922);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n4175, CK => CLK, Q => 
                           n_1373, QN => n19923);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n4174, CK => CLK, Q => 
                           n_1374, QN => n19924);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n4173, CK => CLK, Q => 
                           n_1375, QN => n19925);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n4172, CK => CLK, Q => 
                           n_1376, QN => n19926);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n4171, CK => CLK, Q => 
                           n_1377, QN => n19927);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n4170, CK => CLK, Q => 
                           n_1378, QN => n19928);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n4169, CK => CLK, Q => 
                           n_1379, QN => n19929);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n4168, CK => CLK, Q => 
                           n_1380, QN => n19930);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n4167, CK => CLK, Q => 
                           n_1381, QN => n19931);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n4166, CK => CLK, Q => 
                           n_1382, QN => n19932);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n4165, CK => CLK, Q => 
                           n_1383, QN => n19933);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n4164, CK => CLK, Q => 
                           n_1384, QN => n19934);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n4163, CK => CLK, Q => 
                           n_1385, QN => n19935);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n4162, CK => CLK, Q => 
                           n_1386, QN => n19936);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n4161, CK => CLK, Q => 
                           n_1387, QN => n19937);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n4160, CK => CLK, Q => 
                           n_1388, QN => n19938);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n4159, CK => CLK, Q => 
                           n_1389, QN => n19939);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n4158, CK => CLK, Q => 
                           n_1390, QN => n19940);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n4157, CK => CLK, Q => 
                           n_1391, QN => n19941);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n4156, CK => CLK, Q => 
                           n_1392, QN => n19942);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n4155, CK => CLK, Q => 
                           n_1393, QN => n19943);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n4154, CK => CLK, Q => 
                           n_1394, QN => n19944);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n4153, CK => CLK, Q => 
                           n_1395, QN => n19945);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n4152, CK => CLK, Q => 
                           n_1396, QN => n19946);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n4151, CK => CLK, Q => 
                           n_1397, QN => n19947);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n4150, CK => CLK, Q => 
                           n_1398, QN => n19948);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n4149, CK => CLK, Q => 
                           n_1399, QN => n19949);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n4148, CK => CLK, Q => 
                           n_1400, QN => n19950);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n4147, CK => CLK, Q => 
                           n_1401, QN => n19951);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n4146, CK => CLK, Q => 
                           n_1402, QN => n19952);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n4145, CK => CLK, Q => 
                           n_1403, QN => n19953);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n4144, CK => CLK, Q => 
                           n_1404, QN => n19954);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n4143, CK => CLK, Q => 
                           n_1405, QN => n19955);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n4142, CK => CLK, Q => 
                           n_1406, QN => n19956);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n4141, CK => CLK, Q => 
                           n_1407, QN => n19957);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n4140, CK => CLK, Q => 
                           n_1408, QN => n19958);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n4139, CK => CLK, Q => 
                           n_1409, QN => n19959);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n4138, CK => CLK, Q => 
                           n_1410, QN => n19960);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n4137, CK => CLK, Q => 
                           n_1411, QN => n19961);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n4136, CK => CLK, Q => 
                           n_1412, QN => n19962);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n4135, CK => CLK, Q => 
                           n_1413, QN => n19963);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n4134, CK => CLK, Q => 
                           n21515, QN => n19964);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n4133, CK => CLK, Q => 
                           n21514, QN => n19965);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n4132, CK => CLK, Q => 
                           n21471, QN => n19966);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n4131, CK => CLK, Q => 
                           n21498, QN => n19967);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n4130, CK => CLK, Q => 
                           n21497, QN => n19968);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n4129, CK => CLK, Q => 
                           n21466, QN => n19969);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n4128, CK => CLK, Q => 
                           n21496, QN => n19970);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n4127, CK => CLK, Q => 
                           n21489, QN => n19971);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n4126, CK => CLK, Q => 
                           n21468, QN => n19972);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n4125, CK => CLK, Q => 
                           n21500, QN => n19973);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n4124, CK => CLK, Q => 
                           n21502, QN => n19974);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n4123, CK => CLK, Q => 
                           n21494, QN => n19975);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n4122, CK => CLK, Q => 
                           n21465, QN => n19976);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n4121, CK => CLK, Q => 
                           n21522, QN => n19977);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n4120, CK => CLK, Q => 
                           n21462, QN => n19978);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n4119, CK => CLK, Q => 
                           n21464, QN => n19979);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n4118, CK => CLK, Q => 
                           n21483, QN => n19980);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n4117, CK => CLK, Q => 
                           n21482, QN => n19981);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n4116, CK => CLK, Q => 
                           n21491, QN => n19982);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n4115, CK => CLK, Q => 
                           n21511, QN => n19983);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n4114, CK => CLK, Q => 
                           n21481, QN => n19984);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n4113, CK => CLK, Q => 
                           n21510, QN => n19985);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n4112, CK => CLK, Q => 
                           n21461, QN => n19986);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n4111, CK => CLK, Q => 
                           n21493, QN => n19987);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n4110, CK => CLK, Q => 
                           n21519, QN => n19988);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n4109, CK => CLK, Q => 
                           n21509, QN => n19989);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n4108, CK => CLK, Q => 
                           n21485, QN => n19990);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n4107, CK => CLK, Q => 
                           n21516, QN => n19991);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n4106, CK => CLK, Q => 
                           n21508, QN => n19992);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n4105, CK => CLK, Q => 
                           n21473, QN => n19993);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n4104, CK => CLK, Q => 
                           n21475, QN => n19994);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n4103, CK => CLK, Q => 
                           n21460, QN => n19995);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n4102, CK => CLK, Q => 
                           n21763, QN => n19996);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n4101, CK => CLK, Q => 
                           n21490, QN => n19997);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n4100, CK => CLK, Q => 
                           n21479, QN => n19998);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n4099, CK => CLK, Q => 
                           n21480, QN => n19999);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n4098, CK => CLK, Q => 
                           n21506, QN => n20000);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n4097, CK => CLK, Q => 
                           n21492, QN => n20001);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n4096, CK => CLK, Q => 
                           n21477, QN => n20002);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n4095, CK => CLK, Q => 
                           n21486, QN => n20003);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n4094, CK => CLK, Q => 
                           n21487, QN => n20004);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n4093, CK => CLK, Q => 
                           n21476, QN => n20005);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n4092, CK => CLK, Q => 
                           n21488, QN => n20006);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n4091, CK => CLK, Q => 
                           n21517, QN => n20007);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n4090, CK => CLK, Q => 
                           n21472, QN => n20008);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n4089, CK => CLK, Q => 
                           n21474, QN => n20009);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n4088, CK => CLK, Q => 
                           n21507, QN => n20010);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n4087, CK => CLK, Q => 
                           n21478, QN => n20011);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n4086, CK => CLK, Q => 
                           n21520, QN => n20012);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n4085, CK => CLK, Q => 
                           n21495, QN => n20013);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n4084, CK => CLK, Q => 
                           n21521, QN => n20014);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n4083, CK => CLK, Q => 
                           n21484, QN => n20015);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n4082, CK => CLK, Q => 
                           n21518, QN => n20016);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n4081, CK => CLK, Q => 
                           n21469, QN => n20017);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n4080, CK => CLK, Q => 
                           n21467, QN => n20018);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n4079, CK => CLK, Q => 
                           n21503, QN => n20019);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n4078, CK => CLK, Q => 
                           n21504, QN => n20020);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n4077, CK => CLK, Q => 
                           n21470, QN => n20021);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n4076, CK => CLK, Q => 
                           n21505, QN => n20022);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n4075, CK => CLK, Q => 
                           n21499, QN => n20023);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n4074, CK => CLK, Q => 
                           n21463, QN => n20024);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n4073, CK => CLK, Q => 
                           n21501, QN => n20025);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n4072, CK => CLK, Q => 
                           n21513, QN => n20026);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n4071, CK => CLK, Q => 
                           n21512, QN => n20027);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n4070, CK => CLK, Q => 
                           n20890, QN => n20028);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n4069, CK => CLK, Q => 
                           n20889, QN => n20029);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n4068, CK => CLK, Q => 
                           n20846, QN => n20030);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n4067, CK => CLK, Q => 
                           n20873, QN => n20031);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n4066, CK => CLK, Q => 
                           n20872, QN => n20032);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n4065, CK => CLK, Q => 
                           n20841, QN => n20033);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n4064, CK => CLK, Q => 
                           n20871, QN => n20034);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n4063, CK => CLK, Q => 
                           n20864, QN => n20035);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n4062, CK => CLK, Q => 
                           n20843, QN => n20036);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n4061, CK => CLK, Q => 
                           n20875, QN => n20037);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n4060, CK => CLK, Q => 
                           n20877, QN => n20038);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n4059, CK => CLK, Q => 
                           n20869, QN => n20039);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n4058, CK => CLK, Q => 
                           n20840, QN => n20040);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n4057, CK => CLK, Q => 
                           n20897, QN => n20041);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n4056, CK => CLK, Q => 
                           n20837, QN => n20042);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n4055, CK => CLK, Q => 
                           n20839, QN => n20043);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n4054, CK => CLK, Q => 
                           n20858, QN => n20044);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n4053, CK => CLK, Q => 
                           n20857, QN => n20045);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n4052, CK => CLK, Q => 
                           n20866, QN => n20046);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n4051, CK => CLK, Q => 
                           n20886, QN => n20047);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n4050, CK => CLK, Q => 
                           n20856, QN => n20048);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n4049, CK => CLK, Q => 
                           n20885, QN => n20049);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n4048, CK => CLK, Q => 
                           n20836, QN => n20050);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n4047, CK => CLK, Q => 
                           n20868, QN => n20051);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n4046, CK => CLK, Q => 
                           n20894, QN => n20052);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n4045, CK => CLK, Q => 
                           n20884, QN => n20053);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n4044, CK => CLK, Q => 
                           n20860, QN => n20054);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n4043, CK => CLK, Q => 
                           n20891, QN => n20055);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n4042, CK => CLK, Q => 
                           n20883, QN => n20056);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n4041, CK => CLK, Q => 
                           n20848, QN => n20057);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n4040, CK => CLK, Q => 
                           n20850, QN => n20058);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n4039, CK => CLK, Q => 
                           n20835, QN => n20059);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n4038, CK => CLK, Q => 
                           n20898, QN => n20060);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n4037, CK => CLK, Q => 
                           n20865, QN => n20061);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n4036, CK => CLK, Q => 
                           n20854, QN => n20062);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n4035, CK => CLK, Q => 
                           n20855, QN => n20063);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n4034, CK => CLK, Q => 
                           n20881, QN => n20064);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n4033, CK => CLK, Q => 
                           n20867, QN => n20065);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n4032, CK => CLK, Q => 
                           n20852, QN => n20066);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n4031, CK => CLK, Q => 
                           n20861, QN => n20067);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n4030, CK => CLK, Q => 
                           n20862, QN => n20068);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n4029, CK => CLK, Q => 
                           n20851, QN => n20069);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n4028, CK => CLK, Q => 
                           n20863, QN => n20070);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n4027, CK => CLK, Q => 
                           n20892, QN => n20071);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n4026, CK => CLK, Q => 
                           n20847, QN => n20072);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n4025, CK => CLK, Q => 
                           n20849, QN => n20073);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n4024, CK => CLK, Q => 
                           n20882, QN => n20074);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n4023, CK => CLK, Q => 
                           n20853, QN => n20075);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n4022, CK => CLK, Q => 
                           n20895, QN => n20076);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n4021, CK => CLK, Q => 
                           n20870, QN => n20077);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n4020, CK => CLK, Q => 
                           n20896, QN => n20078);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n4019, CK => CLK, Q => 
                           n20859, QN => n20079);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n4018, CK => CLK, Q => 
                           n20893, QN => n20080);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n4017, CK => CLK, Q => 
                           n20844, QN => n20081);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n4016, CK => CLK, Q => 
                           n20842, QN => n20082);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n4015, CK => CLK, Q => 
                           n20878, QN => n20083);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n4014, CK => CLK, Q => 
                           n20879, QN => n20084);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n4013, CK => CLK, Q => 
                           n20845, QN => n20085);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n4012, CK => CLK, Q => 
                           n20880, QN => n20086);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n4011, CK => CLK, Q => 
                           n20874, QN => n20087);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n4010, CK => CLK, Q => 
                           n20838, QN => n20088);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n4009, CK => CLK, Q => 
                           n20876, QN => n20089);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n4008, CK => CLK, Q => 
                           n20888, QN => n20090);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n4007, CK => CLK, Q => 
                           n20887, QN => n20091);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n4006, CK => CLK, Q => 
                           n21086, QN => n20092);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n4005, CK => CLK, Q => 
                           n21085, QN => n20093);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n4004, CK => CLK, Q => 
                           n21042, QN => n20094);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n4003, CK => CLK, Q => 
                           n21069, QN => n20095);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n4002, CK => CLK, Q => 
                           n21068, QN => n20096);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n4001, CK => CLK, Q => 
                           n21037, QN => n20097);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n4000, CK => CLK, Q => 
                           n21067, QN => n20098);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n3999, CK => CLK, Q => 
                           n21060, QN => n20099);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n3998, CK => CLK, Q => 
                           n21039, QN => n20100);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n3997, CK => CLK, Q => 
                           n21071, QN => n20101);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n3996, CK => CLK, Q => 
                           n21073, QN => n20102);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n3995, CK => CLK, Q => 
                           n21065, QN => n20103);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n3994, CK => CLK, Q => 
                           n21036, QN => n20104);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n3993, CK => CLK, Q => 
                           n21093, QN => n20105);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n3992, CK => CLK, Q => 
                           n21033, QN => n20106);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n3991, CK => CLK, Q => 
                           n21035, QN => n20107);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n3990, CK => CLK, Q => 
                           n21054, QN => n20108);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n3989, CK => CLK, Q => 
                           n21053, QN => n20109);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n3988, CK => CLK, Q => 
                           n21062, QN => n20110);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n3987, CK => CLK, Q => 
                           n21082, QN => n20111);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n3986, CK => CLK, Q => 
                           n21052, QN => n20112);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n3985, CK => CLK, Q => 
                           n21081, QN => n20113);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n3984, CK => CLK, Q => 
                           n21032, QN => n20114);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n3983, CK => CLK, Q => 
                           n21064, QN => n20115);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n3982, CK => CLK, Q => 
                           n21090, QN => n20116);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n3981, CK => CLK, Q => 
                           n21080, QN => n20117);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n3980, CK => CLK, Q => 
                           n21056, QN => n20118);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n3979, CK => CLK, Q => 
                           n21087, QN => n20119);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n3978, CK => CLK, Q => 
                           n21079, QN => n20120);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n3977, CK => CLK, Q => 
                           n21044, QN => n20121);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n3976, CK => CLK, Q => 
                           n21046, QN => n20122);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n3975, CK => CLK, Q => 
                           n21031, QN => n20123);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n3974, CK => CLK, Q => 
                           n21272, QN => n20124);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n3973, CK => CLK, Q => 
                           n21061, QN => n20125);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n3972, CK => CLK, Q => 
                           n21050, QN => n20126);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n3971, CK => CLK, Q => 
                           n21051, QN => n20127);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n3970, CK => CLK, Q => 
                           n21077, QN => n20128);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n3969, CK => CLK, Q => 
                           n21063, QN => n20129);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n3968, CK => CLK, Q => 
                           n21048, QN => n20130);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n3967, CK => CLK, Q => 
                           n21057, QN => n20131);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n3966, CK => CLK, Q => 
                           n21058, QN => n20132);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n3965, CK => CLK, Q => 
                           n21047, QN => n20133);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n3964, CK => CLK, Q => 
                           n21059, QN => n20134);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n3963, CK => CLK, Q => 
                           n21088, QN => n20135);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n3962, CK => CLK, Q => 
                           n21043, QN => n20136);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n3961, CK => CLK, Q => 
                           n21045, QN => n20137);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n3960, CK => CLK, Q => 
                           n21078, QN => n20138);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n3959, CK => CLK, Q => 
                           n21049, QN => n20139);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n3958, CK => CLK, Q => 
                           n21091, QN => n20140);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n3957, CK => CLK, Q => 
                           n21066, QN => n20141);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n3956, CK => CLK, Q => 
                           n21092, QN => n20142);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n3955, CK => CLK, Q => 
                           n21055, QN => n20143);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n3954, CK => CLK, Q => 
                           n21089, QN => n20144);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n3953, CK => CLK, Q => 
                           n21040, QN => n20145);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n3952, CK => CLK, Q => 
                           n21038, QN => n20146);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n3951, CK => CLK, Q => 
                           n21074, QN => n20147);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n3950, CK => CLK, Q => 
                           n21075, QN => n20148);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n3949, CK => CLK, Q => 
                           n21041, QN => n20149);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n3948, CK => CLK, Q => 
                           n21076, QN => n20150);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n3947, CK => CLK, Q => 
                           n21070, QN => n20151);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n3946, CK => CLK, Q => 
                           n21034, QN => n20152);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n3945, CK => CLK, Q => 
                           n21072, QN => n20153);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n3944, CK => CLK, Q => 
                           n21084, QN => n20154);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n3943, CK => CLK, Q => 
                           n21083, QN => n20155);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n3942, CK => CLK, Q => 
                           n_1414, QN => n20156);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n3941, CK => CLK, Q => 
                           n_1415, QN => n20157);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n3940, CK => CLK, Q => 
                           n_1416, QN => n20158);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n3939, CK => CLK, Q => 
                           n_1417, QN => n20159);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n3938, CK => CLK, Q => 
                           n_1418, QN => n20160);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n3937, CK => CLK, Q => 
                           n_1419, QN => n20161);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n3936, CK => CLK, Q => 
                           n_1420, QN => n20162);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n3935, CK => CLK, Q => 
                           n_1421, QN => n20163);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n3934, CK => CLK, Q => 
                           n_1422, QN => n20164);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n3933, CK => CLK, Q => 
                           n_1423, QN => n20165);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n3932, CK => CLK, Q => 
                           n_1424, QN => n20166);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n3931, CK => CLK, Q => 
                           n_1425, QN => n20167);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n3930, CK => CLK, Q => 
                           n_1426, QN => n20168);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n3929, CK => CLK, Q => 
                           n_1427, QN => n20169);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n3928, CK => CLK, Q => 
                           n_1428, QN => n20170);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n3927, CK => CLK, Q => 
                           n_1429, QN => n20171);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n3926, CK => CLK, Q => 
                           n_1430, QN => n20172);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n3925, CK => CLK, Q => 
                           n_1431, QN => n20173);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n3924, CK => CLK, Q => 
                           n_1432, QN => n20174);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n3923, CK => CLK, Q => 
                           n_1433, QN => n20175);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n3922, CK => CLK, Q => 
                           n_1434, QN => n20176);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n3921, CK => CLK, Q => 
                           n_1435, QN => n20177);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n3920, CK => CLK, Q => 
                           n_1436, QN => n20178);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n3919, CK => CLK, Q => 
                           n_1437, QN => n20179);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n3918, CK => CLK, Q => 
                           n_1438, QN => n20180);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n3917, CK => CLK, Q => 
                           n_1439, QN => n20181);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n3916, CK => CLK, Q => 
                           n_1440, QN => n20182);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n3915, CK => CLK, Q => 
                           n_1441, QN => n20183);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n3914, CK => CLK, Q => 
                           n_1442, QN => n20184);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n3913, CK => CLK, Q => 
                           n_1443, QN => n20185);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n3912, CK => CLK, Q => 
                           n_1444, QN => n20186);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n3911, CK => CLK, Q => 
                           n_1445, QN => n20187);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n3910, CK => CLK, Q => 
                           n_1446, QN => n20188);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n3909, CK => CLK, Q => 
                           n_1447, QN => n20189);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n3908, CK => CLK, Q => 
                           n_1448, QN => n20190);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n3907, CK => CLK, Q => 
                           n_1449, QN => n20191);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n3906, CK => CLK, Q => 
                           n_1450, QN => n20192);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n3905, CK => CLK, Q => 
                           n_1451, QN => n20193);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n3904, CK => CLK, Q => 
                           n_1452, QN => n20194);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n3903, CK => CLK, Q => 
                           n_1453, QN => n20195);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n3902, CK => CLK, Q => 
                           n_1454, QN => n20196);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n3901, CK => CLK, Q => 
                           n_1455, QN => n20197);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n3900, CK => CLK, Q => 
                           n_1456, QN => n20198);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n3899, CK => CLK, Q => 
                           n_1457, QN => n20199);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n3898, CK => CLK, Q => 
                           n_1458, QN => n20200);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n3897, CK => CLK, Q => 
                           n_1459, QN => n20201);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n3896, CK => CLK, Q => 
                           n_1460, QN => n20202);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n3895, CK => CLK, Q => 
                           n_1461, QN => n20203);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n3894, CK => CLK, Q => 
                           n_1462, QN => n20204);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n3893, CK => CLK, Q => 
                           n_1463, QN => n20205);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n3892, CK => CLK, Q => 
                           n_1464, QN => n20206);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n3891, CK => CLK, Q => 
                           n_1465, QN => n20207);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n3890, CK => CLK, Q => 
                           n_1466, QN => n20208);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n3889, CK => CLK, Q => 
                           n_1467, QN => n20209);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n3888, CK => CLK, Q => 
                           n_1468, QN => n20210);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n3887, CK => CLK, Q => 
                           n_1469, QN => n20211);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n3886, CK => CLK, Q => 
                           n_1470, QN => n20212);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n3885, CK => CLK, Q => 
                           n_1471, QN => n20213);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n3884, CK => CLK, Q => 
                           n_1472, QN => n20214);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n3883, CK => CLK, Q => 
                           n_1473, QN => n20215);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n3882, CK => CLK, Q => 
                           n_1474, QN => n20216);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n3881, CK => CLK, Q => 
                           n_1475, QN => n20217);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n3880, CK => CLK, Q => 
                           n_1476, QN => n20218);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n3879, CK => CLK, Q => 
                           n_1477, QN => n20219);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n3878, CK => CLK, Q => 
                           n_1478, QN => n20220);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n3877, CK => CLK, Q => 
                           n_1479, QN => n20221);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n3876, CK => CLK, Q => 
                           n_1480, QN => n20222);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n3875, CK => CLK, Q => 
                           n_1481, QN => n20223);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n3874, CK => CLK, Q => 
                           n_1482, QN => n20224);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n3873, CK => CLK, Q => 
                           n_1483, QN => n20225);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n3872, CK => CLK, Q => 
                           n_1484, QN => n20226);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n3871, CK => CLK, Q => 
                           n_1485, QN => n20227);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n3870, CK => CLK, Q => 
                           n_1486, QN => n20228);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n3869, CK => CLK, Q => 
                           n_1487, QN => n20229);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n3868, CK => CLK, Q => 
                           n_1488, QN => n20230);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n3867, CK => CLK, Q => 
                           n_1489, QN => n20231);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n3866, CK => CLK, Q => 
                           n_1490, QN => n20232);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n3865, CK => CLK, Q => 
                           n_1491, QN => n20233);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n3864, CK => CLK, Q => 
                           n_1492, QN => n20234);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n3863, CK => CLK, Q => 
                           n_1493, QN => n20235);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n3862, CK => CLK, Q => 
                           n_1494, QN => n20236);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n3861, CK => CLK, Q => 
                           n_1495, QN => n20237);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n3860, CK => CLK, Q => 
                           n_1496, QN => n20238);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n3859, CK => CLK, Q => 
                           n_1497, QN => n20239);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n3858, CK => CLK, Q => 
                           n_1498, QN => n20240);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n3857, CK => CLK, Q => 
                           n_1499, QN => n20241);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n3856, CK => CLK, Q => 
                           n_1500, QN => n20242);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n3855, CK => CLK, Q => 
                           n_1501, QN => n20243);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n3854, CK => CLK, Q => 
                           n_1502, QN => n20244);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n3853, CK => CLK, Q => 
                           n_1503, QN => n20245);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n3852, CK => CLK, Q => 
                           n_1504, QN => n20246);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n3851, CK => CLK, Q => 
                           n_1505, QN => n20247);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n3850, CK => CLK, Q => 
                           n_1506, QN => n20248);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n3849, CK => CLK, Q => 
                           n_1507, QN => n20249);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n3848, CK => CLK, Q => 
                           n_1508, QN => n20250);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n3847, CK => CLK, Q => 
                           n_1509, QN => n20251);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n3846, CK => CLK, Q => 
                           n_1510, QN => n20252);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n3845, CK => CLK, Q => 
                           n_1511, QN => n20253);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n3844, CK => CLK, Q => 
                           n_1512, QN => n20254);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n3843, CK => CLK, Q => 
                           n_1513, QN => n20255);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n3842, CK => CLK, Q => 
                           n_1514, QN => n20256);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n3841, CK => CLK, Q => 
                           n_1515, QN => n20257);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n3840, CK => CLK, Q => 
                           n_1516, QN => n20258);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n3839, CK => CLK, Q => 
                           n_1517, QN => n20259);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n3838, CK => CLK, Q => 
                           n_1518, QN => n20260);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n3837, CK => CLK, Q => 
                           n_1519, QN => n20261);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n3836, CK => CLK, Q => 
                           n_1520, QN => n20262);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n3835, CK => CLK, Q => 
                           n_1521, QN => n20263);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n3834, CK => CLK, Q => 
                           n_1522, QN => n20264);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n3833, CK => CLK, Q => 
                           n_1523, QN => n20265);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n3832, CK => CLK, Q => 
                           n_1524, QN => n20266);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n3831, CK => CLK, Q => 
                           n_1525, QN => n20267);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n3830, CK => CLK, Q => 
                           n_1526, QN => n20268);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n3829, CK => CLK, Q => 
                           n_1527, QN => n20269);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n3828, CK => CLK, Q => 
                           n_1528, QN => n20270);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n3827, CK => CLK, Q => 
                           n_1529, QN => n20271);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n3826, CK => CLK, Q => 
                           n_1530, QN => n20272);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n3825, CK => CLK, Q => 
                           n_1531, QN => n20273);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n3824, CK => CLK, Q => 
                           n_1532, QN => n20274);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n3823, CK => CLK, Q => 
                           n_1533, QN => n20275);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n3822, CK => CLK, Q => 
                           n_1534, QN => n20276);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n3821, CK => CLK, Q => 
                           n_1535, QN => n20277);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n3820, CK => CLK, Q => 
                           n_1536, QN => n20278);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n3819, CK => CLK, Q => 
                           n_1537, QN => n20279);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n3818, CK => CLK, Q => 
                           n_1538, QN => n20280);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n3817, CK => CLK, Q => 
                           n_1539, QN => n20281);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n3816, CK => CLK, Q => 
                           n_1540, QN => n20282);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n3815, CK => CLK, Q => 
                           n_1541, QN => n20283);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n3814, CK => CLK, Q => 
                           n21899, QN => n20284);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n3813, CK => CLK, Q => 
                           n21898, QN => n20285);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n3812, CK => CLK, Q => 
                           n21858, QN => n20286);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n3811, CK => CLK, Q => 
                           n21895, QN => n20287);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n3810, CK => CLK, Q => 
                           n21894, QN => n20288);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n3809, CK => CLK, Q => 
                           n21856, QN => n20289);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n3808, CK => CLK, Q => 
                           n21891, QN => n20290);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n3807, CK => CLK, Q => 
                           n21875, QN => n20291);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n3806, CK => CLK, Q => 
                           n21854, QN => n20292);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n3805, CK => CLK, Q => 
                           n21888, QN => n20293);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n3804, CK => CLK, Q => 
                           n21887, QN => n20294);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n3803, CK => CLK, Q => 
                           n21886, QN => n20295);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n3802, CK => CLK, Q => 
                           n21851, QN => n20296);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n3801, CK => CLK, Q => 
                           n21906, QN => n20297);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n3800, CK => CLK, Q => 
                           n21850, QN => n20298);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n3799, CK => CLK, Q => 
                           n21849, QN => n20299);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n3798, CK => CLK, Q => 
                           n21873, QN => n20300);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n3797, CK => CLK, Q => 
                           n21871, QN => n20301);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n3796, CK => CLK, Q => 
                           n21870, QN => n20302);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n3795, CK => CLK, Q => 
                           n21883, QN => n20303);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n3794, CK => CLK, Q => 
                           n21869, QN => n20304);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n3793, CK => CLK, Q => 
                           n21882, QN => n20305);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n3792, CK => CLK, Q => 
                           n21846, QN => n20306);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n3791, CK => CLK, Q => 
                           n21881, QN => n20307);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n3790, CK => CLK, Q => 
                           n21902, QN => n20308);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n3789, CK => CLK, Q => 
                           n21880, QN => n20309);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n3788, CK => CLK, Q => 
                           n21863, QN => n20310);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n3787, CK => CLK, Q => 
                           n21900, QN => n20311);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n3786, CK => CLK, Q => 
                           n21877, QN => n20312);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n3785, CK => CLK, Q => 
                           n21845, QN => n20313);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n3784, CK => CLK, Q => 
                           n21860, QN => n20314);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n3783, CK => CLK, Q => 
                           n21844, QN => n20315);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n3782, CK => CLK, Q => 
                           n21907, QN => n20316);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n3781, CK => CLK, Q => 
                           n21859, QN => n20317);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n3780, CK => CLK, Q => 
                           n21861, QN => n20318);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n3779, CK => CLK, Q => 
                           n21862, QN => n20319);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n3778, CK => CLK, Q => 
                           n21878, QN => n20320);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n3777, CK => CLK, Q => 
                           n21879, QN => n20321);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n3776, CK => CLK, Q => 
                           n21864, QN => n20322);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n3775, CK => CLK, Q => 
                           n21865, QN => n20323);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n3774, CK => CLK, Q => 
                           n21866, QN => n20324);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n3773, CK => CLK, Q => 
                           n21867, QN => n20325);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n3772, CK => CLK, Q => 
                           n21868, QN => n20326);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n3771, CK => CLK, Q => 
                           n21901, QN => n20327);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n3770, CK => CLK, Q => 
                           n21847, QN => n20328);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n3769, CK => CLK, Q => 
                           n21848, QN => n20329);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n3768, CK => CLK, Q => 
                           n21884, QN => n20330);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n3767, CK => CLK, Q => 
                           n21872, QN => n20331);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n3766, CK => CLK, Q => 
                           n21904, QN => n20332);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n3765, CK => CLK, Q => 
                           n21885, QN => n20333);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n3764, CK => CLK, Q => 
                           n21905, QN => n20334);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n3763, CK => CLK, Q => 
                           n21874, QN => n20335);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n3762, CK => CLK, Q => 
                           n21903, QN => n20336);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n3761, CK => CLK, Q => 
                           n21852, QN => n20337);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n3760, CK => CLK, Q => 
                           n21853, QN => n20338);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n3759, CK => CLK, Q => 
                           n21889, QN => n20339);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n3758, CK => CLK, Q => 
                           n21890, QN => n20340);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n3757, CK => CLK, Q => 
                           n21855, QN => n20341);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n3756, CK => CLK, Q => 
                           n21892, QN => n20342);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n3755, CK => CLK, Q => 
                           n21893, QN => n20343);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n3754, CK => CLK, Q => 
                           n21857, QN => n20344);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n3753, CK => CLK, Q => 
                           n21896, QN => n20345);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n3752, CK => CLK, Q => 
                           n21897, QN => n20346);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n3751, CK => CLK, Q => 
                           n21876, QN => n20347);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n3750, CK => CLK, Q => 
                           n21018, QN => n20348);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n3749, CK => CLK, Q => 
                           n21017, QN => n20349);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n3748, CK => CLK, Q => 
                           n20977, QN => n20350);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n3747, CK => CLK, Q => 
                           n21014, QN => n20351);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n3746, CK => CLK, Q => 
                           n21013, QN => n20352);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n3745, CK => CLK, Q => 
                           n20975, QN => n20353);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n3744, CK => CLK, Q => 
                           n21010, QN => n20354);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n3743, CK => CLK, Q => 
                           n20994, QN => n20355);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n3742, CK => CLK, Q => 
                           n20973, QN => n20356);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n3741, CK => CLK, Q => 
                           n21007, QN => n20357);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n3740, CK => CLK, Q => 
                           n21006, QN => n20358);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n3739, CK => CLK, Q => 
                           n21005, QN => n20359);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n3738, CK => CLK, Q => 
                           n20970, QN => n20360);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n3737, CK => CLK, Q => 
                           n21025, QN => n20361);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n3736, CK => CLK, Q => 
                           n20969, QN => n20362);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n3735, CK => CLK, Q => 
                           n20968, QN => n20363);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n3734, CK => CLK, Q => 
                           n20992, QN => n20364);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n3733, CK => CLK, Q => 
                           n20990, QN => n20365);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n3732, CK => CLK, Q => 
                           n20989, QN => n20366);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n3731, CK => CLK, Q => 
                           n21002, QN => n20367);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n3730, CK => CLK, Q => 
                           n20988, QN => n20368);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n3729, CK => CLK, Q => 
                           n21001, QN => n20369);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n3728, CK => CLK, Q => 
                           n20965, QN => n20370);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n3727, CK => CLK, Q => 
                           n21000, QN => n20371);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n3726, CK => CLK, Q => 
                           n21021, QN => n20372);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n3725, CK => CLK, Q => 
                           n20999, QN => n20373);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n3724, CK => CLK, Q => 
                           n20982, QN => n20374);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n3723, CK => CLK, Q => 
                           n21019, QN => n20375);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n3722, CK => CLK, Q => 
                           n20996, QN => n20376);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n3721, CK => CLK, Q => 
                           n20964, QN => n20377);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n3720, CK => CLK, Q => 
                           n20979, QN => n20378);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n3719, CK => CLK, Q => 
                           n20963, QN => n20379);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n3718, CK => CLK, Q => 
                           n21026, QN => n20380);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n3717, CK => CLK, Q => 
                           n20978, QN => n20381);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n3716, CK => CLK, Q => 
                           n20980, QN => n20382);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n3715, CK => CLK, Q => 
                           n20981, QN => n20383);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n3714, CK => CLK, Q => 
                           n20997, QN => n20384);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n3713, CK => CLK, Q => 
                           n20998, QN => n20385);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n3712, CK => CLK, Q => 
                           n20983, QN => n20386);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n3711, CK => CLK, Q => 
                           n20984, QN => n20387);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n3710, CK => CLK, Q => 
                           n20985, QN => n20388);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n3709, CK => CLK, Q => 
                           n20986, QN => n20389);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n3708, CK => CLK, Q => 
                           n20987, QN => n20390);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n3707, CK => CLK, Q => 
                           n21020, QN => n20391);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n3706, CK => CLK, Q => 
                           n20966, QN => n20392);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n3705, CK => CLK, Q => 
                           n20967, QN => n20393);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n3704, CK => CLK, Q => 
                           n21003, QN => n20394);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n3703, CK => CLK, Q => 
                           n20991, QN => n20395);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n3702, CK => CLK, Q => 
                           n21023, QN => n20396);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n3701, CK => CLK, Q => 
                           n21004, QN => n20397);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n3700, CK => CLK, Q => 
                           n21024, QN => n20398);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n3699, CK => CLK, Q => 
                           n20993, QN => n20399);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n3698, CK => CLK, Q => 
                           n21022, QN => n20400);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n3697, CK => CLK, Q => 
                           n20971, QN => n20401);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n3696, CK => CLK, Q => 
                           n20972, QN => n20402);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n3695, CK => CLK, Q => 
                           n21008, QN => n20403);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n3694, CK => CLK, Q => 
                           n21009, QN => n20404);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n3693, CK => CLK, Q => 
                           n20974, QN => n20405);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n3692, CK => CLK, Q => 
                           n21011, QN => n20406);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n3691, CK => CLK, Q => 
                           n21012, QN => n20407);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n3690, CK => CLK, Q => 
                           n20976, QN => n20408);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n3689, CK => CLK, Q => 
                           n21015, QN => n20409);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n3688, CK => CLK, Q => 
                           n21016, QN => n20410);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n3687, CK => CLK, Q => 
                           n20995, QN => n20411);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n3686, CK => CLK, Q => 
                           n21352, QN => n20412);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n3685, CK => CLK, Q => 
                           n21354, QN => n20413);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n3684, CK => CLK, Q => 
                           n21356, QN => n20414);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n3683, CK => CLK, Q => 
                           n21358, QN => n20415);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n3682, CK => CLK, Q => 
                           n21360, QN => n20416);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n3681, CK => CLK, Q => 
                           n21362, QN => n20417);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n3680, CK => CLK, Q => 
                           n21364, QN => n20418);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n3679, CK => CLK, Q => 
                           n21366, QN => n20419);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n3678, CK => CLK, Q => 
                           n21368, QN => n20420);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n3677, CK => CLK, Q => 
                           n21370, QN => n20421);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n3676, CK => CLK, Q => 
                           n21372, QN => n20422);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n3675, CK => CLK, Q => 
                           n21374, QN => n20423);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n3674, CK => CLK, Q => 
                           n21376, QN => n20424);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n3673, CK => CLK, Q => 
                           n21378, QN => n20425);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n3672, CK => CLK, Q => 
                           n21380, QN => n20426);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n3671, CK => CLK, Q => 
                           n21382, QN => n20427);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n3670, CK => CLK, Q => 
                           n21384, QN => n20428);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n3669, CK => CLK, Q => 
                           n21386, QN => n20429);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n3668, CK => CLK, Q => 
                           n21388, QN => n20430);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n3667, CK => CLK, Q => 
                           n21390, QN => n20431);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n3666, CK => CLK, Q => 
                           n21392, QN => n20432);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n3665, CK => CLK, Q => 
                           n21394, QN => n20433);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n3664, CK => CLK, Q => 
                           n21396, QN => n20434);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n3663, CK => CLK, Q => 
                           n21398, QN => n20435);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n3662, CK => CLK, Q => 
                           n21400, QN => n20436);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n3661, CK => CLK, Q => 
                           n21402, QN => n20437);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n3660, CK => CLK, Q => 
                           n21404, QN => n20438);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n3659, CK => CLK, Q => 
                           n21406, QN => n20439);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n3658, CK => CLK, Q => 
                           n21408, QN => n20440);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n3657, CK => CLK, Q => 
                           n21410, QN => n20441);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n3656, CK => CLK, Q => 
                           n21412, QN => n20442);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n3655, CK => CLK, Q => 
                           n21414, QN => n20443);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n3654, CK => CLK, Q => 
                           n21351, QN => n20444);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n3653, CK => CLK, Q => 
                           n21413, QN => n20445);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n3652, CK => CLK, Q => 
                           n21411, QN => n20446);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n3651, CK => CLK, Q => 
                           n21409, QN => n20447);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n3650, CK => CLK, Q => 
                           n21407, QN => n20448);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n3649, CK => CLK, Q => 
                           n21405, QN => n20449);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n3648, CK => CLK, Q => 
                           n21403, QN => n20450);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n3647, CK => CLK, Q => 
                           n21401, QN => n20451);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n3646, CK => CLK, Q => 
                           n21399, QN => n20452);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n3645, CK => CLK, Q => 
                           n21397, QN => n20453);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n3644, CK => CLK, Q => 
                           n21395, QN => n20454);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n3643, CK => CLK, Q => 
                           n21393, QN => n20455);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n3642, CK => CLK, Q => 
                           n21391, QN => n20456);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n3641, CK => CLK, Q => 
                           n21389, QN => n20457);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n3640, CK => CLK, Q => 
                           n21387, QN => n20458);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n3639, CK => CLK, Q => 
                           n21385, QN => n20459);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n3638, CK => CLK, Q => 
                           n21383, QN => n20460);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n3637, CK => CLK, Q => 
                           n21381, QN => n20461);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n3636, CK => CLK, Q => 
                           n21379, QN => n20462);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n3635, CK => CLK, Q => 
                           n21377, QN => n20463);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n3634, CK => CLK, Q => 
                           n21375, QN => n20464);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n3633, CK => CLK, Q => 
                           n21373, QN => n20465);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n3632, CK => CLK, Q => 
                           n21371, QN => n20466);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n3631, CK => CLK, Q => 
                           n21369, QN => n20467);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n3630, CK => CLK, Q => 
                           n21367, QN => n20468);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n3629, CK => CLK, Q => 
                           n21365, QN => n20469);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n3628, CK => CLK, Q => 
                           n21363, QN => n20470);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n3627, CK => CLK, Q => 
                           n21361, QN => n20471);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n3626, CK => CLK, Q => 
                           n21359, QN => n20472);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n3625, CK => CLK, Q => 
                           n21357, QN => n20473);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n3624, CK => CLK, Q => 
                           n21355, QN => n20474);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n3623, CK => CLK, Q => 
                           n21353, QN => n20475);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n3622, CK => CLK, Q => 
                           n21973, QN => n20476);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n3621, CK => CLK, Q => 
                           n21975, QN => n20477);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n3620, CK => CLK, Q => 
                           n21977, QN => n20478);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n3619, CK => CLK, Q => 
                           n21979, QN => n20479);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n3618, CK => CLK, Q => 
                           n21981, QN => n20480);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n3617, CK => CLK, Q => 
                           n21983, QN => n20481);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n3616, CK => CLK, Q => 
                           n21985, QN => n20482);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n3615, CK => CLK, Q => 
                           n21987, QN => n20483);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n3614, CK => CLK, Q => 
                           n21989, QN => n20484);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           n21991, QN => n20485);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           n21993, QN => n20486);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           n21995, QN => n20487);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           n21997, QN => n20488);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           n21999, QN => n20489);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           n22001, QN => n20490);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           n22003, QN => n20491);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           n22005, QN => n20492);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           n22007, QN => n20493);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           n22009, QN => n20494);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           n22011, QN => n20495);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           n22013, QN => n20496);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           n22015, QN => n20497);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => 
                           n22017, QN => n20498);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => 
                           n22019, QN => n20499);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => 
                           n22021, QN => n20500);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => 
                           n22023, QN => n20501);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => 
                           n22025, QN => n20502);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => 
                           n22027, QN => n20503);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => 
                           n22029, QN => n20504);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => 
                           n22031, QN => n20505);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => 
                           n22033, QN => n20506);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => 
                           n22035, QN => n20507);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => 
                           n21972, QN => n20508);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => 
                           n22034, QN => n20509);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => 
                           n22032, QN => n20510);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => 
                           n22030, QN => n20511);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => 
                           n22028, QN => n20512);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => 
                           n22026, QN => n20513);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => 
                           n22024, QN => n20514);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => 
                           n22022, QN => n20515);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => 
                           n22020, QN => n20516);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           n22018, QN => n20517);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           n22016, QN => n20518);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           n22014, QN => n20519);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           n22012, QN => n20520);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           n22010, QN => n20521);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           n22008, QN => n20522);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           n22006, QN => n20523);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           n22004, QN => n20524);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           n22002, QN => n20525);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           n22000, QN => n20526);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           n21998, QN => n20527);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           n21996, QN => n20528);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           n21994, QN => n20529);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => 
                           n21992, QN => n20530);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => 
                           n21990, QN => n20531);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => 
                           n21988, QN => n20532);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => 
                           n21986, QN => n20533);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => 
                           n21984, QN => n20534);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => 
                           n21982, QN => n20535);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => 
                           n21980, QN => n20536);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => 
                           n21978, QN => n20537);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => 
                           n21976, QN => n20538);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => 
                           n21974, QN => n20539);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => 
                           n21909, QN => n20540);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => 
                           n21911, QN => n20541);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => 
                           n21913, QN => n20542);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => 
                           n21915, QN => n20543);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => 
                           n21917, QN => n20544);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => 
                           n21919, QN => n20545);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => 
                           n21921, QN => n20546);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => 
                           n21923, QN => n20547);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => 
                           n21925, QN => n20548);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => 
                           n21927, QN => n20549);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => 
                           n21929, QN => n20550);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => 
                           n21931, QN => n20551);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => 
                           n21933, QN => n20552);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => 
                           n21935, QN => n20553);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => 
                           n21937, QN => n20554);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => 
                           n21939, QN => n20555);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => 
                           n21941, QN => n20556);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => 
                           n21943, QN => n20557);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => 
                           n21945, QN => n20558);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => 
                           n21947, QN => n20559);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => 
                           n21949, QN => n20560);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => 
                           n21951, QN => n20561);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => 
                           n21953, QN => n20562);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => 
                           n21955, QN => n20563);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => 
                           n21957, QN => n20564);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => 
                           n21959, QN => n20565);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => 
                           n21961, QN => n20566);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => 
                           n21963, QN => n20567);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => 
                           n21965, QN => n20568);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => 
                           n21967, QN => n20569);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => 
                           n21969, QN => n20570);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => 
                           n21971, QN => n20571);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => 
                           n21908, QN => n20572);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => 
                           n21970, QN => n20573);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => 
                           n21968, QN => n20574);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => 
                           n21966, QN => n20575);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => 
                           n21964, QN => n20576);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => 
                           n21962, QN => n20577);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => 
                           n21960, QN => n20578);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => 
                           n21958, QN => n20579);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => 
                           n21956, QN => n20580);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => 
                           n21954, QN => n20581);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => 
                           n21952, QN => n20582);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => 
                           n21950, QN => n20583);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => 
                           n21948, QN => n20584);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => 
                           n21946, QN => n20585);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => 
                           n21944, QN => n20586);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => 
                           n21942, QN => n20587);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => 
                           n21940, QN => n20588);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => 
                           n21938, QN => n20589);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => 
                           n21936, QN => n20590);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => 
                           n21934, QN => n20591);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => 
                           n21932, QN => n20592);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => 
                           n21930, QN => n20593);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => 
                           n21928, QN => n20594);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => 
                           n21926, QN => n20595);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => 
                           n21924, QN => n20596);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => 
                           n21922, QN => n20597);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => 
                           n21920, QN => n20598);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => 
                           n21918, QN => n20599);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => 
                           n21916, QN => n20600);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => 
                           n21914, QN => n20601);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => 
                           n21912, QN => n20602);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => 
                           n21910, QN => n20603);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => 
                           n20825, QN => n20604);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => 
                           n20824, QN => n20605);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => 
                           n20784, QN => n20606);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => 
                           n20821, QN => n20607);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => 
                           n20820, QN => n20608);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => 
                           n20782, QN => n20609);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => 
                           n20817, QN => n20610);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => 
                           n20801, QN => n20611);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => 
                           n20780, QN => n20612);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => 
                           n20814, QN => n20613);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => 
                           n20813, QN => n20614);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => 
                           n20812, QN => n20615);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => 
                           n20777, QN => n20616);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => 
                           n20832, QN => n20617);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => 
                           n20776, QN => n20618);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => 
                           n20775, QN => n20619);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => 
                           n20799, QN => n20620);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => 
                           n20797, QN => n20621);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => 
                           n20796, QN => n20622);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => 
                           n20809, QN => n20623);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => 
                           n20795, QN => n20624);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => 
                           n20808, QN => n20625);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => 
                           n20772, QN => n20626);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => 
                           n20807, QN => n20627);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => 
                           n20828, QN => n20628);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => 
                           n20806, QN => n20629);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => 
                           n20789, QN => n20630);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => 
                           n20826, QN => n20631);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => 
                           n20803, QN => n20632);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => 
                           n20771, QN => n20633);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => 
                           n20786, QN => n20634);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => 
                           n20770, QN => n20635);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => 
                           n20833, QN => n20636);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => 
                           n20785, QN => n20637);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => 
                           n20787, QN => n20638);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => 
                           n20788, QN => n20639);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => 
                           n20804, QN => n20640);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => 
                           n20805, QN => n20641);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => 
                           n20790, QN => n20642);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => 
                           n20791, QN => n20643);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => 
                           n20792, QN => n20644);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => 
                           n20793, QN => n20645);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => 
                           n20794, QN => n20646);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => 
                           n20827, QN => n20647);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => 
                           n20773, QN => n20648);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => 
                           n20774, QN => n20649);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => 
                           n20810, QN => n20650);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => 
                           n20798, QN => n20651);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => 
                           n20830, QN => n20652);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => 
                           n20811, QN => n20653);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => 
                           n20831, QN => n20654);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => 
                           n20800, QN => n20655);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => 
                           n20829, QN => n20656);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => 
                           n20778, QN => n20657);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => 
                           n20779, QN => n20658);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => 
                           n20815, QN => n20659);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => 
                           n20816, QN => n20660);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => 
                           n20781, QN => n20661);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => 
                           n20818, QN => n20662);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => 
                           n20819, QN => n20663);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => 
                           n20783, QN => n20664);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => 
                           n20822, QN => n20665);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => 
                           n20823, QN => n20666);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => 
                           n20802, QN => n20667);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => 
                           n21342, QN => n20668);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => 
                           n21341, QN => n20669);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => 
                           n21301, QN => n20670);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => 
                           n21338, QN => n20671);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => 
                           n21337, QN => n20672);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => 
                           n21299, QN => n20673);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => 
                           n21334, QN => n20674);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => 
                           n21318, QN => n20675);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => 
                           n21297, QN => n20676);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => 
                           n21331, QN => n20677);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => 
                           n21330, QN => n20678);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => 
                           n21329, QN => n20679);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => 
                           n21294, QN => n20680);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => 
                           n21349, QN => n20681);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => 
                           n21293, QN => n20682);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => 
                           n21292, QN => n20683);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => 
                           n21316, QN => n20684);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => 
                           n21314, QN => n20685);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => 
                           n21313, QN => n20686);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => 
                           n21326, QN => n20687);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => 
                           n21312, QN => n20688);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => 
                           n21325, QN => n20689);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => 
                           n21289, QN => n20690);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => 
                           n21324, QN => n20691);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => 
                           n21345, QN => n20692);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => 
                           n21323, QN => n20693);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => 
                           n21306, QN => n20694);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => 
                           n21343, QN => n20695);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => 
                           n21320, QN => n20696);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => 
                           n21288, QN => n20697);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => 
                           n21303, QN => n20698);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => 
                           n21287, QN => n20699);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => 
                           n21350, QN => n20700);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => 
                           n21302, QN => n20701);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => 
                           n21304, QN => n20702);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => 
                           n21305, QN => n20703);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => 
                           n21321, QN => n20704);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => 
                           n21322, QN => n20705);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => 
                           n21307, QN => n20706);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => 
                           n21308, QN => n20707);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => 
                           n21309, QN => n20708);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => 
                           n21310, QN => n20709);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => 
                           n21311, QN => n20710);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => 
                           n21344, QN => n20711);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => 
                           n21290, QN => n20712);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => 
                           n21291, QN => n20713);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => 
                           n21327, QN => n20714);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => 
                           n21315, QN => n20715);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => 
                           n21347, QN => n20716);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => 
                           n21328, QN => n20717);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => 
                           n21348, QN => n20718);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => 
                           n21317, QN => n20719);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => 
                           n21346, QN => n20720);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => 
                           n21295, QN => n20721);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => 
                           n21296, QN => n20722);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => 
                           n21332, QN => n20723);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => 
                           n21333, QN => n20724);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => 
                           n21298, QN => n20725);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => 
                           n21335, QN => n20726);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => 
                           n21336, QN => n20727);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => 
                           n21300, QN => n20728);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => 
                           n21339, QN => n20729);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => 
                           n21340, QN => n20730);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => 
                           n21319, QN => n20731);
   CWP_reg_4_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => CWP_4_port, QN
                           => n994);
   CWP_reg_5_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => CWP_5_port, QN
                           => n993);
   CWP_reg_6_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => CWP_6_port, QN
                           => n992);
   CWP_reg_7_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => CWP_7_port, QN
                           => n991);
   CWP_reg_8_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => CWP_8_port, QN
                           => n990);
   CWP_reg_9_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => CWP_9_port, QN
                           => n989);
   CWP_reg_10_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => CWP_10_port, 
                           QN => n988);
   CWP_reg_11_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => CWP_11_port, 
                           QN => n987);
   CWP_reg_12_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => CWP_12_port, 
                           QN => n986);
   CWP_reg_13_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => CWP_13_port, 
                           QN => n985);
   CWP_reg_14_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => CWP_14_port, 
                           QN => n984);
   CWP_reg_15_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => CWP_15_port, 
                           QN => n983);
   CWP_reg_16_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => CWP_16_port, 
                           QN => n982);
   CWP_reg_17_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => CWP_17_port, 
                           QN => n981);
   CWP_reg_18_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => CWP_18_port, 
                           QN => n980);
   CWP_reg_19_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => CWP_19_port, 
                           QN => n979);
   CWP_reg_20_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => CWP_20_port, 
                           QN => n978);
   CWP_reg_21_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => CWP_21_port, 
                           QN => n977);
   CWP_reg_22_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => CWP_22_port, 
                           QN => n976);
   CWP_reg_23_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => CWP_23_port, 
                           QN => n975);
   CWP_reg_24_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => CWP_24_port, 
                           QN => n974);
   CWP_reg_25_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => CWP_25_port, 
                           QN => n973);
   CWP_reg_26_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => CWP_26_port, 
                           QN => n972);
   CWP_reg_27_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => CWP_27_port, 
                           QN => n971);
   CWP_reg_28_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => CWP_28_port, 
                           QN => n970);
   CWP_reg_29_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => CWP_29_port, 
                           QN => n969);
   CWP_reg_30_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => CWP_30_port, 
                           QN => n968);
   CWP_reg_31_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => CWP_31_port, 
                           QN => n967);
   n13243 <= '0';
   n13244 <= '1';
   n13245 <= '0';
   n13246 <= '0';
   n13247 <= '0';
   n13248 <= '1';
   U11075 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => n25409, A3 => n25407, ZN
                           => n15181);
   U11076 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n25408, A3 => n25407, ZN
                           => n15180);
   U11080 : NAND3_X1 port map( A1 => n23945, A2 => n23284, A3 => n16579, ZN => 
                           n16529);
   r286 : REGISTER_FILE_WINDOWING_DW01_addsub_0 port map( A(31) => i_31_port, 
                           A(30) => i_30_port, A(29) => i_29_port, A(28) => 
                           i_28_port, A(27) => i_27_port, A(26) => i_26_port, 
                           A(25) => i_25_port, A(24) => i_24_port, A(23) => 
                           i_23_port, A(22) => i_22_port, A(21) => i_21_port, 
                           A(20) => i_20_port, A(19) => i_19_port, A(18) => 
                           i_18_port, A(17) => i_17_port, A(16) => i_16_port, 
                           A(15) => i_15_port, A(14) => i_14_port, A(13) => 
                           i_13_port, A(12) => i_12_port, A(11) => i_11_port, 
                           A(10) => i_10_port, A(9) => i_9_port, A(8) => 
                           i_8_port, A(7) => i_7_port, A(6) => i_6_port, A(5) 
                           => i_5_port, A(4) => i_4_port, A(3) => i_3_port, 
                           A(2) => n24143, A(1) => i_1_port, A(0) => i_0_port, 
                           B(31) => n13243, B(30) => n13243, B(29) => n13243, 
                           B(28) => n13243, B(27) => n13243, B(26) => n13243, 
                           B(25) => n13243, B(24) => n13243, B(23) => n13243, 
                           B(22) => n13243, B(21) => n13243, B(20) => n13243, 
                           B(19) => n13243, B(18) => n13243, B(17) => n13243, 
                           B(16) => n13243, B(15) => n13243, B(14) => n13243, 
                           B(13) => n13243, B(12) => n13243, B(11) => n13243, 
                           B(10) => n13243, B(9) => n13243, B(8) => n13243, 
                           B(7) => n13243, B(6) => n13243, B(5) => n13243, B(4)
                           => n13243, B(3) => n13243, B(2) => n13243, B(1) => 
                           n13243, B(0) => n13244, CI => n13247, ADD_SUB => 
                           n13247, SUM(31) => N653, SUM(30) => N652, SUM(29) =>
                           N651, SUM(28) => N650, SUM(27) => N649, SUM(26) => 
                           N648, SUM(25) => N647, SUM(24) => N646, SUM(23) => 
                           N645, SUM(22) => N644, SUM(21) => N643, SUM(20) => 
                           N642, SUM(19) => N641, SUM(18) => N640, SUM(17) => 
                           N639, SUM(16) => N638, SUM(15) => N637, SUM(14) => 
                           N636, SUM(13) => N635, SUM(12) => N634, SUM(11) => 
                           N633, SUM(10) => N632, SUM(9) => N631, SUM(8) => 
                           N630, SUM(7) => N629, SUM(6) => N628, SUM(5) => N627
                           , SUM(4) => N626, SUM(3) => N625, SUM(2) => N624, 
                           SUM(1) => N623, SUM(0) => n_1542, CO => n_1543);
   r268 : REGISTER_FILE_WINDOWING_DW01_cmp6_0 port map( A(31) => U3_U2_Z_31, 
                           A(30) => U3_U2_Z_30, A(29) => U3_U2_Z_29, A(28) => 
                           U3_U2_Z_28, A(27) => U3_U2_Z_27, A(26) => U3_U2_Z_26
                           , A(25) => U3_U2_Z_25, A(24) => U3_U2_Z_24, A(23) =>
                           U3_U2_Z_23, A(22) => U3_U2_Z_22, A(21) => U3_U2_Z_21
                           , A(20) => U3_U2_Z_20, A(19) => U3_U2_Z_19, A(18) =>
                           U3_U2_Z_18, A(17) => U3_U2_Z_17, A(16) => U3_U2_Z_16
                           , A(15) => U3_U2_Z_15, A(14) => U3_U2_Z_14, A(13) =>
                           U3_U2_Z_13, A(12) => U3_U2_Z_12, A(11) => U3_U2_Z_11
                           , A(10) => U3_U2_Z_10, A(9) => U3_U2_Z_9, A(8) => 
                           U3_U2_Z_8, A(7) => U3_U2_Z_7, A(6) => U3_U2_Z_6, 
                           A(5) => U3_U2_Z_5, A(4) => U3_U2_Z_4, A(3) => 
                           U3_U2_Z_3, A(2) => U3_U2_Z_2, A(1) => U3_U2_Z_1, 
                           A(0) => U3_U2_Z_0, B(31) => U3_U3_Z_31, B(30) => 
                           U3_U3_Z_30, B(29) => U3_U3_Z_29, B(28) => U3_U3_Z_28
                           , B(27) => U3_U3_Z_27, B(26) => U3_U3_Z_26, B(25) =>
                           U3_U3_Z_25, B(24) => U3_U3_Z_24, B(23) => U3_U3_Z_23
                           , B(22) => U3_U3_Z_22, B(21) => U3_U3_Z_21, B(20) =>
                           U3_U3_Z_20, B(19) => U3_U3_Z_19, B(18) => U3_U3_Z_18
                           , B(17) => U3_U3_Z_17, B(16) => U3_U3_Z_16, B(15) =>
                           U3_U3_Z_15, B(14) => U3_U3_Z_14, B(13) => U3_U3_Z_13
                           , B(12) => U3_U3_Z_12, B(11) => U3_U3_Z_11, B(10) =>
                           U3_U3_Z_10, B(9) => U3_U3_Z_9, B(8) => U3_U3_Z_8, 
                           B(7) => U3_U3_Z_7, B(6) => U3_U3_Z_6, B(5) => 
                           U3_U3_Z_5, B(4) => U3_U3_Z_4, B(3) => U3_U3_Z_3, 
                           B(2) => U3_U3_Z_2, B(1) => U3_U3_Z_1, B(0) => 
                           U3_U3_Z_0, TC => n13248, LT => N2739, GT => n_1544, 
                           EQ => N139, LE => n_1545, GE => n_1546, NE => n_1547
                           );
   r235 : REGISTER_FILE_WINDOWING_DW01_addsub_2 port map( A(31) => U3_U7_Z_31, 
                           A(30) => U3_U7_Z_30, A(29) => U3_U7_Z_29, A(28) => 
                           U3_U7_Z_28, A(27) => U3_U7_Z_27, A(26) => U3_U7_Z_26
                           , A(25) => U3_U7_Z_25, A(24) => U3_U7_Z_24, A(23) =>
                           U3_U7_Z_23, A(22) => U3_U7_Z_22, A(21) => U3_U7_Z_21
                           , A(20) => U3_U7_Z_20, A(19) => U3_U7_Z_19, A(18) =>
                           U3_U7_Z_18, A(17) => U3_U7_Z_17, A(16) => U3_U7_Z_16
                           , A(15) => U3_U7_Z_15, A(14) => U3_U7_Z_14, A(13) =>
                           U3_U7_Z_13, A(12) => U3_U7_Z_12, A(11) => U3_U7_Z_11
                           , A(10) => U3_U7_Z_10, A(9) => U3_U7_Z_9, A(8) => 
                           U3_U7_Z_8, A(7) => U3_U7_Z_7, A(6) => U3_U7_Z_6, 
                           A(5) => U3_U7_Z_5, A(4) => U3_U7_Z_4, A(3) => 
                           U3_U7_Z_3, A(2) => U3_U7_Z_2, A(1) => U3_U7_Z_1, 
                           A(0) => U3_U7_Z_0, B(31) => n13243, B(30) => n13243,
                           B(29) => n13243, B(28) => n13243, B(27) => n13243, 
                           B(26) => n13243, B(25) => n13243, B(24) => n13243, 
                           B(23) => n13243, B(22) => n13243, B(21) => n13243, 
                           B(20) => n13243, B(19) => n13243, B(18) => n13243, 
                           B(17) => n13243, B(16) => n13243, B(15) => n13243, 
                           B(14) => n13243, B(13) => n13243, B(12) => n13243, 
                           B(11) => n13243, B(10) => n13243, B(9) => n13243, 
                           B(8) => n13243, B(7) => n13243, B(6) => n13243, B(5)
                           => n13243, B(4) => n13243, B(3) => U3_U8_Z_3, B(2) 
                           => U3_U8_Z_2, B(1) => n20764, B(0) => U3_U8_Z_0, CI 
                           => n13246, ADD_SUB => U3_U9_Z_0, SUM(31) => N241, 
                           SUM(30) => N240, SUM(29) => N239, SUM(28) => N238, 
                           SUM(27) => N237, SUM(26) => N236, SUM(25) => N235, 
                           SUM(24) => N234, SUM(23) => N233, SUM(22) => N232, 
                           SUM(21) => N231, SUM(20) => N230, SUM(19) => N229, 
                           SUM(18) => N228, SUM(17) => N227, SUM(16) => N226, 
                           SUM(15) => N225, SUM(14) => N224, SUM(13) => N223, 
                           SUM(12) => N222, SUM(11) => N221, SUM(10) => N220, 
                           SUM(9) => N219, SUM(8) => N218, SUM(7) => N217, 
                           SUM(6) => N216, SUM(5) => N215, SUM(4) => N214, 
                           SUM(3) => N213, SUM(2) => N212, SUM(1) => N211, 
                           SUM(0) => N210, CO => n_1548);
   r233 : REGISTER_FILE_WINDOWING_DW01_add_0 port map( A(31) => CWP_31_port, 
                           A(30) => CWP_30_port, A(29) => CWP_29_port, A(28) =>
                           CWP_28_port, A(27) => CWP_27_port, A(26) => 
                           CWP_26_port, A(25) => CWP_25_port, A(24) => 
                           CWP_24_port, A(23) => CWP_23_port, A(22) => 
                           CWP_22_port, A(21) => CWP_21_port, A(20) => 
                           CWP_20_port, A(19) => CWP_19_port, A(18) => 
                           CWP_18_port, A(17) => CWP_17_port, A(16) => 
                           CWP_16_port, A(15) => CWP_15_port, A(14) => 
                           CWP_14_port, A(13) => CWP_13_port, A(12) => 
                           CWP_12_port, A(11) => CWP_11_port, A(10) => 
                           CWP_10_port, A(9) => CWP_9_port, A(8) => CWP_8_port,
                           A(7) => CWP_7_port, A(6) => CWP_6_port, A(5) => 
                           CWP_5_port, A(4) => CWP_4_port, A(3) => CWP_3_port, 
                           A(2) => CWP_2_port, A(1) => CWP_1_port, A(0) => 
                           CWP_0_port, B(31) => U3_U1_Z_31, B(30) => U3_U1_Z_30
                           , B(29) => U3_U1_Z_29, B(28) => U3_U1_Z_28, B(27) =>
                           U3_U1_Z_27, B(26) => U3_U1_Z_26, B(25) => U3_U1_Z_25
                           , B(24) => U3_U1_Z_24, B(23) => U3_U1_Z_23, B(22) =>
                           U3_U1_Z_22, B(21) => U3_U1_Z_21, B(20) => U3_U1_Z_20
                           , B(19) => U3_U1_Z_19, B(18) => U3_U1_Z_18, B(17) =>
                           U3_U1_Z_17, B(16) => U3_U1_Z_16, B(15) => U3_U1_Z_15
                           , B(14) => U3_U1_Z_14, B(13) => U3_U1_Z_13, B(12) =>
                           U3_U1_Z_12, B(11) => U3_U1_Z_11, B(10) => U3_U1_Z_10
                           , B(9) => U3_U1_Z_9, B(8) => U3_U1_Z_8, B(7) => 
                           U3_U1_Z_7, B(6) => U3_U1_Z_6, B(5) => U3_U1_Z_5, 
                           B(4) => U3_U1_Z_4, B(3) => U3_U1_Z_3, B(2) => 
                           U3_U1_Z_2, B(1) => U3_U1_Z_1, B(0) => U3_U1_Z_0, CI 
                           => n13245, SUM(31) => N106, SUM(30) => N105, SUM(29)
                           => N104, SUM(28) => N103, SUM(27) => N102, SUM(26) 
                           => N101, SUM(25) => N100, SUM(24) => N99, SUM(23) =>
                           N98, SUM(22) => N97, SUM(21) => N96, SUM(20) => N95,
                           SUM(19) => N94, SUM(18) => N93, SUM(17) => N92, 
                           SUM(16) => N91, SUM(15) => N90, SUM(14) => N89, 
                           SUM(13) => N88, SUM(12) => N87, SUM(11) => N86, 
                           SUM(10) => N85, SUM(9) => N84, SUM(8) => N83, SUM(7)
                           => N82, SUM(6) => N81, SUM(5) => N80, SUM(4) => N79,
                           SUM(3) => N78, SUM(2) => N77, SUM(1) => N76, SUM(0) 
                           => N75, CO => n_1549);
   CWP_reg_0_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => CWP_0_port, QN
                           => n3046);
   i_reg_8_inst : DFF_X1 port map( D => n13234, CK => CLK, Q => i_8_port, QN =>
                           n3256);
   i_reg_9_inst : DFF_X1 port map( D => n13233, CK => CLK, Q => i_9_port, QN =>
                           n3255);
   i_reg_19_inst : DFF_X1 port map( D => n13223, CK => CLK, Q => i_19_port, QN 
                           => n3271);
   i_reg_20_inst : DFF_X1 port map( D => n13222, CK => CLK, Q => i_20_port, QN 
                           => n3270);
   i_reg_21_inst : DFF_X1 port map( D => n13221, CK => CLK, Q => i_21_port, QN 
                           => n3269);
   i_reg_1_inst : DFF_X1 port map( D => n13241, CK => CLK, Q => i_1_port, QN =>
                           n22673);
   i_reg_4_inst : DFF_X1 port map( D => n13238, CK => CLK, Q => i_4_port, QN =>
                           n3252);
   FILLING_reg : DFF_X1 port map( D => n5641, CK => CLK, Q => n24003, QN => 
                           n5700);
   SWP_reg_16_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => n_1550, QN =>
                           n22780);
   SWP_reg_13_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => n22533, QN =>
                           n22781);
   SWP_reg_3_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => n_1551, QN => 
                           n22784);
   SWP_reg_0_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => n_1552, QN => 
                           n22788);
   SWP_reg_1_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => n_1553, QN => 
                           n22982);
   SWP_reg_2_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => n_1554, QN => 
                           n22983);
   SPILLING_reg : DFF_X1 port map( D => n5642, CK => CLK, Q => n20834, QN => 
                           n5699);
   OUT1_reg_37_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => OUT1_37_port
                           , QN => n24965);
   OUT1_reg_0_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1555);
   OUT1_reg_40_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => OUT1_40_port
                           , QN => n25013);
   OUT1_reg_36_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => OUT1_36_port
                           , QN => n24949);
   OUT1_reg_22_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => OUT1_22_port
                           , QN => n24725);
   OUT1_reg_63_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => OUT1_63_port
                           , QN => n25393);
   OUT1_reg_25_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => OUT1_25_port
                           , QN => n24773);
   OUT1_reg_21_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => OUT1_21_port
                           , QN => n24709);
   OUT1_reg_24_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => OUT1_24_port
                           , QN => n24757);
   OUT1_reg_8_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => OUT1_8_port, 
                           QN => n24501);
   OUT1_reg_59_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => OUT1_59_port
                           , QN => n25317);
   OUT1_reg_52_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => OUT1_52_port
                           , QN => n25205);
   OUT1_reg_50_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => OUT1_50_port
                           , QN => n25173);
   OUT1_reg_48_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => OUT1_48_port
                           , QN => n25141);
   OUT1_reg_46_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => OUT1_46_port
                           , QN => n25109);
   OUT1_reg_43_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => OUT1_43_port
                           , QN => n25061);
   OUT1_reg_27_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => OUT1_27_port
                           , QN => n24805);
   OUT1_reg_9_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => OUT1_9_port, 
                           QN => n24517);
   OUT1_reg_2_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => OUT1_2_port, 
                           QN => n24405);
   OUT1_reg_62_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => OUT1_62_port
                           , QN => n25365);
   OUT1_reg_58_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => OUT1_58_port
                           , QN => n25301);
   OUT1_reg_49_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => OUT1_49_port
                           , QN => n25157);
   OUT1_reg_45_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => OUT1_45_port
                           , QN => n25093);
   OUT1_reg_42_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => OUT1_42_port
                           , QN => n25045);
   OUT1_reg_20_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => OUT1_20_port
                           , QN => n24693);
   OUT1_reg_16_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => OUT1_16_port
                           , QN => n24629);
   OUT1_reg_34_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => OUT1_34_port
                           , QN => n24917);
   OUT1_reg_18_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => OUT1_18_port
                           , QN => n24661);
   OUT1_reg_41_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => OUT1_41_port
                           , QN => n25029);
   OUT1_reg_39_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => OUT1_39_port
                           , QN => n24997);
   OUT1_reg_33_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => OUT1_33_port
                           , QN => n24901);
   OUT1_reg_17_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => OUT1_17_port
                           , QN => n24645);
   OUT1_reg_15_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => OUT1_15_port
                           , QN => n24613);
   OUT1_reg_13_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => OUT1_13_port
                           , QN => n24581);
   OUT1_reg_7_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => OUT1_7_port, 
                           QN => n24485);
   OUT1_reg_32_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => OUT1_32_port
                           , QN => n24885);
   OUT1_reg_14_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => OUT1_14_port
                           , QN => n24597);
   OUT1_reg_11_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => OUT1_11_port
                           , QN => n24549);
   OUT1_reg_61_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => OUT1_61_port
                           , QN => n25349);
   OUT1_reg_28_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => OUT1_28_port
                           , QN => n24821);
   OUT1_reg_26_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => OUT1_26_port
                           , QN => n24789);
   OUT1_reg_5_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => OUT1_5_port, 
                           QN => n24453);
   OUT1_reg_60_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => OUT1_60_port
                           , QN => n25333);
   OUT1_reg_54_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => OUT1_54_port
                           , QN => n25237);
   OUT1_reg_47_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => OUT1_47_port
                           , QN => n25125);
   OUT1_reg_38_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => OUT1_38_port
                           , QN => n24981);
   OUT1_reg_31_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => OUT1_31_port
                           , QN => n24869);
   OUT1_reg_29_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => OUT1_29_port
                           , QN => n24837);
   OUT1_reg_23_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => OUT1_23_port
                           , QN => n24741);
   OUT1_reg_6_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => OUT1_6_port, 
                           QN => n24469);
   OUT1_reg_4_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => OUT1_4_port, 
                           QN => n24437);
   OUT1_reg_57_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => OUT1_57_port
                           , QN => n25285);
   OUT1_reg_55_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => OUT1_55_port
                           , QN => n25253);
   OUT1_reg_53_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => OUT1_53_port
                           , QN => n25221);
   OUT1_reg_51_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => OUT1_51_port
                           , QN => n25189);
   OUT1_reg_44_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => OUT1_44_port
                           , QN => n25077);
   OUT1_reg_30_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => OUT1_30_port
                           , QN => n24853);
   OUT1_reg_12_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => OUT1_12_port
                           , QN => n24565);
   OUT1_reg_56_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => OUT1_56_port
                           , QN => n25269);
   OUT1_reg_35_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => OUT1_35_port
                           , QN => n24933);
   OUT1_reg_10_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => OUT1_10_port
                           , QN => n24533);
   OUT1_reg_19_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => OUT1_19_port
                           , QN => n24677);
   OUT1_reg_3_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => OUT1_3_port, 
                           QN => n24421);
   OUT1_reg_1_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => OUT1_1_port, 
                           QN => n24389);
   SWP_reg_15_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => n20756, QN =>
                           n24065);
   CWP_reg_3_inst : DFF_X2 port map( D => n5415, CK => CLK, Q => CWP_3_port, QN
                           => n3043);
   CWP_reg_2_inst : DFF_X2 port map( D => n5417, CK => CLK, Q => CWP_2_port, QN
                           => n3045);
   SWP_reg_10_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => n20761, QN =>
                           n24073);
   SWP_reg_12_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => n20759, QN =>
                           n24069);
   SWP_reg_17_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => n20754, QN =>
                           n24062);
   SWP_reg_11_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => n20760, QN =>
                           n24071);
   SWP_reg_18_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => n20753, QN =>
                           n24060);
   SWP_reg_19_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => n20752, QN =>
                           n24058);
   SWP_reg_29_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => n_1556, QN =>
                           n24047);
   SWP_reg_30_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => n_1557, QN =>
                           n24045);
   MEM_BUS_reg_4_inst : DFF_X1 port map( D => n22764, CK => CLK, Q => 
                           MEM_BUS_4_port, QN => n_1558);
   MEM_BUS_reg_3_inst : DFF_X1 port map( D => n22763, CK => CLK, Q => 
                           MEM_BUS_3_port, QN => n_1559);
   MEM_BUS_reg_2_inst : DFF_X1 port map( D => n22762, CK => CLK, Q => 
                           MEM_BUS_2_port, QN => n_1560);
   MEM_BUS_reg_1_inst : DFF_X1 port map( D => n22761, CK => CLK, Q => 
                           MEM_BUS_1_port, QN => n_1561);
   MEM_BUS_reg_63_inst : DFF_X1 port map( D => n22759, CK => CLK, Q => 
                           MEM_BUS_63_port, QN => n_1562);
   MEM_BUS_reg_62_inst : DFF_X1 port map( D => n22758, CK => CLK, Q => 
                           MEM_BUS_62_port, QN => n_1563);
   MEM_BUS_reg_61_inst : DFF_X1 port map( D => n22757, CK => CLK, Q => 
                           MEM_BUS_61_port, QN => n_1564);
   MEM_BUS_reg_60_inst : DFF_X1 port map( D => n22756, CK => CLK, Q => 
                           MEM_BUS_60_port, QN => n_1565);
   MEM_BUS_reg_59_inst : DFF_X1 port map( D => n22755, CK => CLK, Q => 
                           MEM_BUS_59_port, QN => n_1566);
   MEM_BUS_reg_58_inst : DFF_X1 port map( D => n22754, CK => CLK, Q => 
                           MEM_BUS_58_port, QN => n_1567);
   MEM_BUS_reg_57_inst : DFF_X1 port map( D => n22753, CK => CLK, Q => 
                           MEM_BUS_57_port, QN => n_1568);
   MEM_BUS_reg_56_inst : DFF_X1 port map( D => n22752, CK => CLK, Q => 
                           MEM_BUS_56_port, QN => n_1569);
   MEM_BUS_reg_55_inst : DFF_X1 port map( D => n22751, CK => CLK, Q => 
                           MEM_BUS_55_port, QN => n_1570);
   MEM_BUS_reg_54_inst : DFF_X1 port map( D => n22750, CK => CLK, Q => 
                           MEM_BUS_54_port, QN => n_1571);
   MEM_BUS_reg_53_inst : DFF_X1 port map( D => n22749, CK => CLK, Q => 
                           MEM_BUS_53_port, QN => n_1572);
   MEM_BUS_reg_52_inst : DFF_X1 port map( D => n22748, CK => CLK, Q => 
                           MEM_BUS_52_port, QN => n_1573);
   MEM_BUS_reg_51_inst : DFF_X1 port map( D => n22747, CK => CLK, Q => 
                           MEM_BUS_51_port, QN => n_1574);
   MEM_BUS_reg_50_inst : DFF_X1 port map( D => n22746, CK => CLK, Q => 
                           MEM_BUS_50_port, QN => n_1575);
   MEM_BUS_reg_49_inst : DFF_X1 port map( D => n22745, CK => CLK, Q => 
                           MEM_BUS_49_port, QN => n_1576);
   MEM_BUS_reg_48_inst : DFF_X1 port map( D => n22744, CK => CLK, Q => 
                           MEM_BUS_48_port, QN => n_1577);
   MEM_BUS_reg_47_inst : DFF_X1 port map( D => n22743, CK => CLK, Q => 
                           MEM_BUS_47_port, QN => n_1578);
   MEM_BUS_reg_46_inst : DFF_X1 port map( D => n22742, CK => CLK, Q => 
                           MEM_BUS_46_port, QN => n_1579);
   MEM_BUS_reg_45_inst : DFF_X1 port map( D => n22741, CK => CLK, Q => 
                           MEM_BUS_45_port, QN => n_1580);
   MEM_BUS_reg_44_inst : DFF_X1 port map( D => n22740, CK => CLK, Q => 
                           MEM_BUS_44_port, QN => n_1581);
   MEM_BUS_reg_43_inst : DFF_X1 port map( D => n22739, CK => CLK, Q => 
                           MEM_BUS_43_port, QN => n_1582);
   MEM_BUS_reg_42_inst : DFF_X1 port map( D => n22738, CK => CLK, Q => 
                           MEM_BUS_42_port, QN => n_1583);
   MEM_BUS_reg_41_inst : DFF_X1 port map( D => n22737, CK => CLK, Q => 
                           MEM_BUS_41_port, QN => n_1584);
   MEM_BUS_reg_40_inst : DFF_X1 port map( D => n22736, CK => CLK, Q => 
                           MEM_BUS_40_port, QN => n_1585);
   MEM_BUS_reg_39_inst : DFF_X1 port map( D => n22735, CK => CLK, Q => 
                           MEM_BUS_39_port, QN => n_1586);
   MEM_BUS_reg_38_inst : DFF_X1 port map( D => n22734, CK => CLK, Q => 
                           MEM_BUS_38_port, QN => n_1587);
   MEM_BUS_reg_37_inst : DFF_X1 port map( D => n22733, CK => CLK, Q => 
                           MEM_BUS_37_port, QN => n_1588);
   MEM_BUS_reg_36_inst : DFF_X1 port map( D => n22732, CK => CLK, Q => 
                           MEM_BUS_36_port, QN => n_1589);
   MEM_BUS_reg_35_inst : DFF_X1 port map( D => n22731, CK => CLK, Q => 
                           MEM_BUS_35_port, QN => n_1590);
   MEM_BUS_reg_34_inst : DFF_X1 port map( D => n22730, CK => CLK, Q => 
                           MEM_BUS_34_port, QN => n_1591);
   MEM_BUS_reg_33_inst : DFF_X1 port map( D => n22729, CK => CLK, Q => 
                           MEM_BUS_33_port, QN => n_1592);
   MEM_BUS_reg_32_inst : DFF_X1 port map( D => n22728, CK => CLK, Q => 
                           MEM_BUS_32_port, QN => n_1593);
   MEM_BUS_reg_31_inst : DFF_X1 port map( D => n22727, CK => CLK, Q => 
                           MEM_BUS_31_port, QN => n_1594);
   MEM_BUS_reg_30_inst : DFF_X1 port map( D => n22726, CK => CLK, Q => 
                           MEM_BUS_30_port, QN => n_1595);
   MEM_BUS_reg_29_inst : DFF_X1 port map( D => n22725, CK => CLK, Q => 
                           MEM_BUS_29_port, QN => n_1596);
   MEM_BUS_reg_28_inst : DFF_X1 port map( D => n22724, CK => CLK, Q => 
                           MEM_BUS_28_port, QN => n_1597);
   MEM_BUS_reg_27_inst : DFF_X1 port map( D => n22723, CK => CLK, Q => 
                           MEM_BUS_27_port, QN => n_1598);
   MEM_BUS_reg_26_inst : DFF_X1 port map( D => n22722, CK => CLK, Q => 
                           MEM_BUS_26_port, QN => n_1599);
   MEM_BUS_reg_25_inst : DFF_X1 port map( D => n22721, CK => CLK, Q => 
                           MEM_BUS_25_port, QN => n_1600);
   MEM_BUS_reg_24_inst : DFF_X1 port map( D => n22720, CK => CLK, Q => 
                           MEM_BUS_24_port, QN => n_1601);
   MEM_BUS_reg_23_inst : DFF_X1 port map( D => n22719, CK => CLK, Q => 
                           MEM_BUS_23_port, QN => n_1602);
   MEM_BUS_reg_22_inst : DFF_X1 port map( D => n22718, CK => CLK, Q => 
                           MEM_BUS_22_port, QN => n_1603);
   MEM_BUS_reg_21_inst : DFF_X1 port map( D => n22717, CK => CLK, Q => 
                           MEM_BUS_21_port, QN => n_1604);
   MEM_BUS_reg_20_inst : DFF_X1 port map( D => n22716, CK => CLK, Q => 
                           MEM_BUS_20_port, QN => n_1605);
   MEM_BUS_reg_19_inst : DFF_X1 port map( D => n22715, CK => CLK, Q => 
                           MEM_BUS_19_port, QN => n_1606);
   MEM_BUS_reg_18_inst : DFF_X1 port map( D => n22714, CK => CLK, Q => 
                           MEM_BUS_18_port, QN => n_1607);
   MEM_BUS_reg_17_inst : DFF_X1 port map( D => n22713, CK => CLK, Q => 
                           MEM_BUS_17_port, QN => n_1608);
   MEM_BUS_reg_16_inst : DFF_X1 port map( D => n22712, CK => CLK, Q => 
                           MEM_BUS_16_port, QN => n_1609);
   MEM_BUS_reg_15_inst : DFF_X1 port map( D => n22711, CK => CLK, Q => 
                           MEM_BUS_15_port, QN => n_1610);
   MEM_BUS_reg_14_inst : DFF_X1 port map( D => n22710, CK => CLK, Q => 
                           MEM_BUS_14_port, QN => n_1611);
   MEM_BUS_reg_13_inst : DFF_X1 port map( D => n22709, CK => CLK, Q => 
                           MEM_BUS_13_port, QN => n_1612);
   MEM_BUS_reg_12_inst : DFF_X1 port map( D => n22708, CK => CLK, Q => 
                           MEM_BUS_12_port, QN => n_1613);
   MEM_BUS_reg_11_inst : DFF_X1 port map( D => n22707, CK => CLK, Q => 
                           MEM_BUS_11_port, QN => n_1614);
   MEM_BUS_reg_10_inst : DFF_X1 port map( D => n22706, CK => CLK, Q => 
                           MEM_BUS_10_port, QN => n_1615);
   MEM_BUS_reg_9_inst : DFF_X1 port map( D => n22705, CK => CLK, Q => 
                           MEM_BUS_9_port, QN => n_1616);
   MEM_BUS_reg_8_inst : DFF_X1 port map( D => n22704, CK => CLK, Q => 
                           MEM_BUS_8_port, QN => n_1617);
   MEM_BUS_reg_7_inst : DFF_X1 port map( D => n22703, CK => CLK, Q => 
                           MEM_BUS_7_port, QN => n_1618);
   U11116 : AND4_X1 port map( A1 => n20765, A2 => n20766, A3 => n20767, A4 => 
                           n20768, ZN => n24005);
   U11117 : AND4_X1 port map( A1 => n969, A2 => n970, A3 => n968, A4 => n967, 
                           ZN => n20765);
   U11118 : AND4_X1 port map( A1 => n973, A2 => n974, A3 => n971, A4 => n972, 
                           ZN => n20766);
   U11119 : AND4_X1 port map( A1 => n977, A2 => n978, A3 => n975, A4 => n976, 
                           ZN => n20767);
   U11120 : AND4_X1 port map( A1 => n981, A2 => n982, A3 => n979, A4 => n980, 
                           ZN => n20768);
   U11121 : BUF_X1 port map( A => N2739, Z => n20769);
   U11122 : AND4_X1 port map( A1 => n3253, A2 => n3242, A3 => n3252, A4 => 
                           n3251, ZN => n22551);
   U11123 : AND4_X1 port map( A1 => n993, A2 => n994, A3 => n991, A4 => n992, 
                           ZN => n22537);
   U11124 : AND4_X1 port map( A1 => n3046, A2 => n3045, A3 => n3043, A4 => 
                           n3044, ZN => n22538);
   U11125 : AND4_X1 port map( A1 => n989, A2 => n990, A3 => n987, A4 => n988, 
                           ZN => n22536);
   U11126 : AND2_X1 port map( A1 => n16552, A2 => n23329, ZN => n15212);
   U11127 : AND2_X1 port map( A1 => n16552, A2 => n23318, ZN => n15211);
   U11128 : AND4_X1 port map( A1 => n22788, A2 => n22794, A3 => n22982, A4 => 
                           n22983, ZN => n22557);
   U11129 : AND4_X1 port map( A1 => n22784, A2 => n22787, A3 => n22791, A4 => 
                           n22792, ZN => n22556);
   U11130 : AND4_X1 port map( A1 => n3268, A2 => n3246, A3 => n3245, A4 => 
                           n3244, ZN => n22526);
   U11131 : AND4_X1 port map( A1 => n3260, A2 => n3267, A3 => n3266, A4 => 
                           n3265, ZN => n22548);
   U11132 : AND4_X1 port map( A1 => n3241, A2 => n3263, A3 => n3262, A4 => 
                           n3261, ZN => n22549);
   U11133 : AND4_X1 port map( A1 => n3258, A2 => n3257, A3 => n3256, A4 => 
                           n3255, ZN => n22550);
   U11134 : AND2_X1 port map( A1 => n23329, A2 => n16555, ZN => n15221);
   U11135 : AND2_X1 port map( A1 => n23318, A2 => n16555, ZN => n15222);
   U11136 : OAI221_X1 port map( B1 => n24090, B2 => n22784, C1 => n3043, C2 => 
                           n23009, A => n24080, ZN => U3_U7_Z_3);
   U11137 : BUF_X2 port map( A => n23014, Z => n23012);
   U11138 : NAND2_X1 port map( A1 => n24091, A2 => n22628, ZN => U3_U9_Z_0);
   U11139 : NAND3_X1 port map( A1 => n24356, A2 => ADD_RD1(0), A3 => n24352, ZN
                           => n25385);
   U11140 : AND2_X1 port map( A1 => n23032, A2 => N221, ZN => U3_U1_Z_11);
   U11141 : AND2_X1 port map( A1 => N217, A2 => n23032, ZN => U3_U1_Z_7);
   U11142 : AND2_X1 port map( A1 => n23032, A2 => N215, ZN => U3_U1_Z_5);
   U11143 : OAI221_X1 port map( B1 => n22770, B2 => n24060, C1 => n980, C2 => 
                           n23008, A => n24059, ZN => U3_U7_Z_18);
   U11144 : OAI221_X1 port map( B1 => n22777, B2 => n22795, C1 => n975, C2 => 
                           n23007, A => n24053, ZN => U3_U7_Z_23);
   U11145 : OAI221_X1 port map( B1 => n22778, B2 => n22793, C1 => n976, C2 => 
                           n23007, A => n24054, ZN => U3_U7_Z_22);
   U11146 : BUF_X1 port map( A => n23055, Z => n23048);
   U11147 : BUF_X1 port map( A => n23046, Z => n23044);
   U11148 : BUF_X1 port map( A => n23055, Z => n23049);
   U11149 : BUF_X1 port map( A => n23046, Z => n23043);
   U11150 : BUF_X1 port map( A => n23055, Z => n23050);
   U11151 : BUF_X1 port map( A => n23047, Z => n23042);
   U11152 : BUF_X1 port map( A => n23054, Z => n23051);
   U11153 : BUF_X1 port map( A => n23047, Z => n23041);
   U11154 : BUF_X1 port map( A => n23054, Z => n23052);
   U11155 : BUF_X1 port map( A => n23047, Z => n23040);
   U11156 : AND4_X1 port map( A1 => n22535, A2 => n22536, A3 => n22537, A4 => 
                           n22538, ZN => n24006);
   U11157 : AND4_X1 port map( A1 => n985, A2 => n986, A3 => n983, A4 => n984, 
                           ZN => n22535);
   U11158 : BUF_X1 port map( A => n24097, Z => n23026);
   U11159 : BUF_X2 port map( A => n22963, Z => n22801);
   U11160 : AOI22_X2 port map( A1 => MEM_BUSread(62), A2 => n23050, B1 => 
                           DATAIN(62), B2 => n23045, ZN => n16664);
   U11161 : AOI22_X2 port map( A1 => MEM_BUSread(60), A2 => n23048, B1 => 
                           DATAIN(60), B2 => n23045, ZN => n16663);
   U11162 : AOI22_X2 port map( A1 => MEM_BUSread(58), A2 => n23048, B1 => 
                           DATAIN(58), B2 => n23045, ZN => n16662);
   U11163 : AOI22_X2 port map( A1 => MEM_BUSread(56), A2 => n23048, B1 => 
                           DATAIN(56), B2 => n23045, ZN => n16661);
   U11164 : AOI22_X2 port map( A1 => MEM_BUSread(54), A2 => n23048, B1 => 
                           DATAIN(54), B2 => n23044, ZN => n16660);
   U11165 : AOI22_X2 port map( A1 => MEM_BUSread(52), A2 => n23048, B1 => 
                           DATAIN(52), B2 => n23044, ZN => n16659);
   U11166 : AOI22_X2 port map( A1 => MEM_BUSread(36), A2 => n23049, B1 => 
                           DATAIN(36), B2 => n23044, ZN => n16651);
   U11167 : AOI22_X2 port map( A1 => MEM_BUSread(34), A2 => n23049, B1 => 
                           DATAIN(34), B2 => n23044, ZN => n16650);
   U11168 : AOI22_X2 port map( A1 => MEM_BUSread(32), A2 => n23049, B1 => 
                           DATAIN(32), B2 => n23044, ZN => n16649);
   U11169 : AOI22_X2 port map( A1 => MEM_BUSread(30), A2 => n23049, B1 => 
                           DATAIN(30), B2 => n23043, ZN => n16648);
   U11170 : AOI22_X2 port map( A1 => MEM_BUSread(28), A2 => n23049, B1 => 
                           DATAIN(28), B2 => n23043, ZN => n16647);
   U11171 : AOI22_X2 port map( A1 => MEM_BUSread(12), A2 => n23050, B1 => 
                           DATAIN(12), B2 => n23043, ZN => n16639);
   U11172 : AOI22_X2 port map( A1 => MEM_BUSread(10), A2 => n23050, B1 => 
                           DATAIN(10), B2 => n23043, ZN => n16638);
   U11173 : AOI22_X2 port map( A1 => MEM_BUSread(8), A2 => n23050, B1 => 
                           DATAIN(8), B2 => n23043, ZN => n16637);
   U11174 : AOI22_X2 port map( A1 => MEM_BUSread(6), A2 => n23050, B1 => 
                           DATAIN(6), B2 => n23042, ZN => n16636);
   U11175 : AOI22_X2 port map( A1 => MEM_BUSread(9), A2 => n23051, B1 => 
                           DATAIN(9), B2 => n23042, ZN => n16628);
   U11176 : AOI22_X2 port map( A1 => MEM_BUSread(11), A2 => n23051, B1 => 
                           DATAIN(11), B2 => n23042, ZN => n16627);
   U11177 : AOI22_X2 port map( A1 => MEM_BUSread(13), A2 => n23051, B1 => 
                           DATAIN(13), B2 => n23042, ZN => n16626);
   U11178 : AOI22_X2 port map( A1 => MEM_BUSread(15), A2 => n23051, B1 => 
                           DATAIN(15), B2 => n23042, ZN => n16625);
   U11179 : AOI22_X2 port map( A1 => MEM_BUSread(17), A2 => n23051, B1 => 
                           DATAIN(17), B2 => n23041, ZN => n16624);
   U11180 : AOI22_X2 port map( A1 => MEM_BUSread(33), A2 => n23052, B1 => 
                           DATAIN(33), B2 => n23041, ZN => n16616);
   U11181 : AOI22_X2 port map( A1 => MEM_BUSread(35), A2 => n23052, B1 => 
                           DATAIN(35), B2 => n23041, ZN => n16615);
   U11182 : AOI22_X2 port map( A1 => MEM_BUSread(37), A2 => n23052, B1 => 
                           DATAIN(37), B2 => n23041, ZN => n16614);
   U11183 : AOI22_X2 port map( A1 => MEM_BUSread(39), A2 => n23052, B1 => 
                           DATAIN(39), B2 => n23041, ZN => n16613);
   U11184 : AOI22_X2 port map( A1 => MEM_BUSread(41), A2 => n23052, B1 => 
                           DATAIN(41), B2 => n23040, ZN => n16612);
   U11185 : AOI22_X2 port map( A1 => MEM_BUSread(57), A2 => n23053, B1 => 
                           DATAIN(57), B2 => n23040, ZN => n16604);
   U11186 : AOI22_X2 port map( A1 => MEM_BUSread(59), A2 => n23053, B1 => 
                           DATAIN(59), B2 => n23040, ZN => n16603);
   U11187 : AOI22_X2 port map( A1 => MEM_BUSread(61), A2 => n23053, B1 => 
                           DATAIN(61), B2 => n23040, ZN => n16602);
   U11188 : AOI22_X2 port map( A1 => MEM_BUSread(63), A2 => n23053, B1 => 
                           DATAIN(63), B2 => n23040, ZN => n16601);
   U11189 : CLKBUF_X3 port map( A => n25381, Z => n22937);
   U11190 : OAI222_X1 port map( A1 => n23024, A2 => n24026, B1 => n24116, B2 =>
                           n23019, C1 => n985, C2 => n23017, ZN => n3357);
   U11191 : BUF_X1 port map( A => n5699, Z => n22768);
   U11192 : AND2_X1 port map( A1 => n24008, A2 => n24003, ZN => n21415);
   U11193 : NAND2_X1 port map( A1 => n23006, A2 => n24085, ZN => n21429);
   U11194 : AND3_X1 port map( A1 => n24331, A2 => n24335, A3 => n24332, ZN => 
                           n21438);
   U11195 : AND3_X1 port map( A1 => n24331, A2 => n24333, A3 => n24332, ZN => 
                           n21440);
   U11196 : AND3_X1 port map( A1 => n24336, A2 => n24335, A3 => n24334, ZN => 
                           n21443);
   U11197 : AND3_X1 port map( A1 => n24336, A2 => n24334, A3 => n24333, ZN => 
                           n21444);
   U11198 : AND2_X1 port map( A1 => n24359, A2 => n24173, ZN => n21445);
   U11199 : AND2_X1 port map( A1 => n24173, A2 => n24361, ZN => n21447);
   U11200 : AND2_X1 port map( A1 => n21447, A2 => n23468, ZN => n21448);
   U11201 : AND2_X1 port map( A1 => n23507, A2 => n21447, ZN => n21450);
   U11202 : AND2_X1 port map( A1 => n23436, A2 => n21447, ZN => n21451);
   U11203 : AND2_X1 port map( A1 => n21447, A2 => n23413, ZN => n21452);
   U11204 : AND2_X1 port map( A1 => n24359, A2 => n24360, ZN => n21454);
   U11205 : AND2_X1 port map( A1 => n23270, A2 => n23283, ZN => n21456);
   U11206 : AND2_X1 port map( A1 => n23285, A2 => n24003, ZN => n21457);
   U11207 : AND2_X1 port map( A1 => n5700, A2 => n23283, ZN => n21458);
   U11208 : AND3_X1 port map( A1 => n24342, A2 => n22690, A3 => n22493, ZN => 
                           n21459);
   U11209 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => n24368, ZN => n22484);
   U11210 : AND2_X1 port map( A1 => n24131, A2 => WR, ZN => n22485);
   U11211 : AND2_X1 port map( A1 => n24355, A2 => n24368, ZN => n22486);
   U11212 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n24369,
                           ZN => n22487);
   U11213 : CLKBUF_X1 port map( A => n23026, Z => n23023);
   U11214 : CLKBUF_X1 port map( A => n23026, Z => n23025);
   U11215 : NOR2_X1 port map( A1 => n24351, A2 => ADD_RD1(1), ZN => n22488);
   U11216 : NOR2_X1 port map( A1 => n24351, A2 => ADD_RD1(1), ZN => n22932);
   U11217 : CLKBUF_X1 port map( A => n22502, Z => n23030);
   U11218 : NAND4_X1 port map( A1 => n24087, A2 => n24008, A3 => n22512, A4 => 
                           n24003, ZN => n24090);
   U11219 : INV_X1 port map( A => n22489, ZN => n24092);
   U11220 : OAI222_X4 port map( A1 => n23025, A2 => n24023, B1 => n22504, B2 =>
                           n23019, C1 => n988, C2 => n23017, ZN => n3360);
   U11221 : AND3_X2 port map( A1 => n22512, A2 => n24002, A3 => n20834, ZN => 
                           n22489);
   U11222 : CLKBUF_X1 port map( A => N77, Z => n22490);
   U11223 : AND2_X1 port map( A1 => n22957, A2 => n21285, ZN => n22491);
   U11224 : AND2_X1 port map( A1 => n23275, A2 => n20962, ZN => n22492);
   U11225 : NOR3_X1 port map( A1 => n22491, A2 => n22492, A3 => n24357, ZN => 
                           n24373);
   U11226 : BUF_X2 port map( A => n22956, Z => n22957);
   U11227 : BUF_X1 port map( A => n23030, Z => n23028);
   U11228 : BUF_X1 port map( A => n23030, Z => n23029);
   U11229 : BUF_X1 port map( A => n24087, Z => n22510);
   U11230 : CLKBUF_X1 port map( A => n24341, Z => n22493);
   U11231 : INV_X2 port map( A => N79, ZN => n24179);
   U11232 : AND3_X4 port map( A1 => n22488, A2 => ADD_RD1(0), A3 => n24369, ZN 
                           => n22494);
   U11233 : AND2_X1 port map( A1 => n23032, A2 => N224, ZN => U3_U1_Z_14);
   U11234 : CLKBUF_X1 port map( A => N214, Z => n22495);
   U11235 : CLKBUF_X1 port map( A => n24090, Z => n23015);
   U11236 : CLKBUF_X1 port map( A => n23015, Z => n22770);
   U11237 : AND4_X1 port map( A1 => n22674, A2 => i_2_port, A3 => n3254, A4 => 
                           n3247, ZN => n22496);
   U11238 : AND4_X1 port map( A1 => i_2_port, A2 => n22674, A3 => n3254, A4 => 
                           n3247, ZN => n22524);
   U11239 : CLKBUF_X3 port map( A => n23014, Z => n23013);
   U11240 : CLKBUF_X1 port map( A => n24184, Z => n22497);
   U11241 : CLKBUF_X1 port map( A => N211, Z => n22498);
   U11242 : AND4_X1 port map( A1 => n22496, A2 => n22525, A3 => n22526, A4 => 
                           n22527, ZN => n22499);
   U11243 : AND4_X1 port map( A1 => n22524, A2 => n22525, A3 => n22526, A4 => 
                           n22527, ZN => n23947);
   U11244 : CLKBUF_X1 port map( A => n24110, Z => n22500);
   U11245 : BUF_X1 port map( A => n23030, Z => n23027);
   U11246 : INV_X1 port map( A => n22502, ZN => n24093);
   U11247 : BUF_X1 port map( A => n22691, Z => n23010);
   U11248 : AND2_X1 port map( A1 => n24356, A2 => n22487, ZN => n22501);
   U11249 : AND3_X1 port map( A1 => n24341, A2 => n24008, A3 => n24003, ZN => 
                           n22502);
   U11250 : CLKBUF_X1 port map( A => N217, Z => n22503);
   U11251 : INV_X1 port map( A => n22528, ZN => n22504);
   U11252 : OAI222_X1 port map( A1 => n23023, A2 => n24041, B1 => n24101, B2 =>
                           n23021, C1 => n970, C2 => n23016, ZN => n3342);
   U11253 : BUF_X2 port map( A => n23282, Z => n23275);
   U11254 : CLKBUF_X1 port map( A => n24185, Z => n22505);
   U11255 : CLKBUF_X1 port map( A => N210, Z => n22506);
   U11256 : AND2_X1 port map( A1 => n24091, A2 => n22628, ZN => n22507);
   U11257 : AND2_X1 port map( A1 => n23032, A2 => N233, ZN => U3_U1_Z_23);
   U11258 : INV_X1 port map( A => n24179, ZN => n22508);
   U11259 : CLKBUF_X3 port map( A => n25389, Z => n22951);
   U11260 : CLKBUF_X3 port map( A => n25381, Z => n22935);
   U11261 : CLKBUF_X3 port map( A => n23014, Z => n23011);
   U11262 : CLKBUF_X1 port map( A => N216, Z => n22511);
   U11263 : AND2_X2 port map( A1 => n23948, A2 => n23947, ZN => n22512);
   U11264 : CLKBUF_X1 port map( A => N225, Z => n22513);
   U11265 : AND2_X1 port map( A1 => n23032, A2 => N213, ZN => U3_U1_Z_3);
   U11266 : CLKBUF_X3 port map( A => n25388, Z => n22964);
   U11267 : CLKBUF_X3 port map( A => n25388, Z => n22966);
   U11268 : CLKBUF_X3 port map( A => n25388, Z => n22967);
   U11269 : CLKBUF_X3 port map( A => n25388, Z => n22965);
   U11270 : OR2_X1 port map( A1 => n24346, A2 => n24347, ZN => n22514);
   U11271 : OR2_X1 port map( A1 => n24346, A2 => n24347, ZN => n22515);
   U11272 : BUF_X2 port map( A => n22514, Z => n22516);
   U11273 : BUF_X2 port map( A => n22514, Z => n22517);
   U11274 : BUF_X2 port map( A => n22515, Z => n22518);
   U11275 : BUF_X2 port map( A => n22515, Z => n22519);
   U11276 : BUF_X2 port map( A => n25378, Z => n22520);
   U11277 : BUF_X2 port map( A => n25378, Z => n22521);
   U11278 : OR2_X1 port map( A1 => n24346, A2 => n24347, ZN => n25378);
   U11279 : BUF_X2 port map( A => n25383, Z => n22522);
   U11280 : BUF_X2 port map( A => n25383, Z => n22523);
   U11281 : AND3_X1 port map( A1 => N2739, A2 => ADD_RD1(3), A3 => n21456, ZN 
                           => n22696);
   U11282 : AND4_X1 port map( A1 => n3243, A2 => n3250, A3 => n3249, A4 => 
                           n3248, ZN => n22525);
   U11283 : AND4_X1 port map( A1 => n3264, A2 => n3271, A3 => n3270, A4 => 
                           n3269, ZN => n22527);
   U11284 : CLKBUF_X1 port map( A => N220, Z => n22528);
   U11285 : INV_X1 port map( A => n23991, ZN => n22529);
   U11286 : CLKBUF_X1 port map( A => N223, Z => n22530);
   U11287 : CLKBUF_X1 port map( A => n24120, Z => n22531);
   U11288 : CLKBUF_X1 port map( A => N212, Z => n22532);
   U11289 : NOR4_X1 port map( A1 => n20754, A2 => n20753, A3 => n20752, A4 => 
                           n20750, ZN => n22554);
   U11290 : NOR4_X1 port map( A1 => n20760, A2 => n20759, A3 => n22533, A4 => 
                           n22534, ZN => n22555);
   U11291 : AND4_X1 port map( A1 => n22554, A2 => n22555, A3 => n22556, A4 => 
                           n22557, ZN => n23990);
   U11292 : AND2_X1 port map( A1 => n23032, A2 => N225, ZN => U3_U1_Z_15);
   U11293 : INV_X1 port map( A => n24124, ZN => n22542);
   U11294 : CLKBUF_X3 port map( A => n25381, Z => n22936);
   U11295 : CLKBUF_X3 port map( A => n25381, Z => n22934);
   U11296 : CLKBUF_X3 port map( A => n25385, Z => n22980);
   U11297 : BUF_X2 port map( A => n25383, Z => n22921);
   U11298 : CLKBUF_X3 port map( A => n25387, Z => n22639);
   U11299 : NAND2_X1 port map( A1 => n22696, A2 => ADD_RD1(0), ZN => n22543);
   U11300 : OR2_X2 port map( A1 => n22543, A2 => n22544, ZN => n25384);
   U11301 : OR2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), ZN => n22544);
   U11302 : NAND4_X1 port map( A1 => WR, A2 => n22700, A3 => n24008, A4 => 
                           n24130, ZN => n22545);
   U11303 : NAND4_X1 port map( A1 => WR, A2 => n22700, A3 => n24008, A4 => 
                           n24130, ZN => n22546);
   U11304 : CLKBUF_X1 port map( A => N213, Z => n22547);
   U11305 : NAND4_X1 port map( A1 => WR, A2 => n22700, A3 => n24008, A4 => 
                           n24130, ZN => n24126);
   U11306 : AND2_X1 port map( A1 => N216, A2 => n23032, ZN => U3_U1_Z_6);
   U11307 : INV_X2 port map( A => n24086, ZN => n24008);
   U11308 : AND4_X2 port map( A1 => n22548, A2 => n22549, A3 => n22550, A4 => 
                           n22551, ZN => n23948);
   U11309 : AND2_X1 port map( A1 => n22916, A2 => n22191, ZN => n22552);
   U11310 : AND2_X1 port map( A1 => n22802, A2 => n21183, ZN => n22553);
   U11311 : NOR3_X1 port map( A1 => n22552, A2 => n22553, A3 => n24435, ZN => 
                           n24441);
   U11312 : OAI222_X1 port map( A1 => n23024, A2 => n24024, B1 => n24118, B2 =>
                           n23019, C1 => n987, C2 => n23017, ZN => n3359);
   U11313 : AND2_X1 port map( A1 => n22922, A2 => n22186, ZN => n22558);
   U11314 : AND2_X1 port map( A1 => n22969, A2 => n21269, ZN => n22559);
   U11315 : NOR3_X1 port map( A1 => n22558, A2 => n22559, A3 => n24882, ZN => 
                           n24890);
   U11316 : AND2_X1 port map( A1 => n22912, A2 => n22202, ZN => n22560);
   U11317 : AND2_X1 port map( A1 => n22804, A2 => n21175, ZN => n22561);
   U11318 : NOR3_X1 port map( A1 => n22560, A2 => n22561, A3 => n24755, ZN => 
                           n24761);
   U11319 : AND2_X1 port map( A1 => n22917, A2 => n22210, ZN => n22562);
   U11320 : AND2_X1 port map( A1 => n22812, A2 => n21177, ZN => n22563);
   U11321 : NOR3_X1 port map( A1 => n22562, A2 => n22563, A3 => n25123, ZN => 
                           n25129);
   U11322 : BUF_X2 port map( A => n22910, Z => n22917);
   U11323 : AND2_X1 port map( A1 => n22914, A2 => n22222, ZN => n22564);
   U11324 : AND2_X1 port map( A1 => n22806, A2 => n21205, ZN => n22565);
   U11325 : NOR3_X1 port map( A1 => n22564, A2 => n22565, A3 => n25347, ZN => 
                           n25353);
   U11326 : AND2_X1 port map( A1 => n22922, A2 => n22189, ZN => n22566);
   U11327 : AND2_X1 port map( A1 => n22969, A2 => n21268, ZN => n22567);
   U11328 : NOR3_X1 port map( A1 => n22566, A2 => n22567, A3 => n25010, ZN => 
                           n25018);
   U11329 : AND2_X1 port map( A1 => n22921, A2 => n22187, ZN => n22568);
   U11330 : AND2_X1 port map( A1 => n22969, A2 => n21270, ZN => n22569);
   U11331 : NOR3_X1 port map( A1 => n22568, A2 => n22569, A3 => n24946, ZN => 
                           n24954);
   U11332 : AND2_X1 port map( A1 => n22522, A2 => n22185, ZN => n22570);
   U11333 : AND2_X1 port map( A1 => n22969, A2 => n21267, ZN => n22571);
   U11334 : NOR3_X1 port map( A1 => n22570, A2 => n22571, A3 => n24610, ZN => 
                           n24618);
   U11335 : AND2_X1 port map( A1 => n22912, A2 => n22223, ZN => n22572);
   U11336 : AND2_X1 port map( A1 => n22805, A2 => n21206, ZN => n22573);
   U11337 : NOR3_X1 port map( A1 => n22572, A2 => n22573, A3 => n25386, ZN => 
                           n25398);
   U11338 : BUF_X1 port map( A => n22910, Z => n22912);
   U11339 : AND2_X1 port map( A1 => n22918, A2 => n22203, ZN => n22574);
   U11340 : AND2_X1 port map( A1 => n22803, A2 => n21195, ZN => n22575);
   U11341 : NOR3_X1 port map( A1 => n22574, A2 => n22575, A3 => n24771, ZN => 
                           n24777);
   U11342 : BUF_X1 port map( A => n22910, Z => n22918);
   U11343 : AND2_X1 port map( A1 => n22914, A2 => n22204, ZN => n22576);
   U11344 : AND2_X1 port map( A1 => n22802, A2 => n21176, ZN => n22577);
   U11345 : NOR3_X1 port map( A1 => n22576, A2 => n22577, A3 => n24787, ZN => 
                           n24793);
   U11346 : BUF_X1 port map( A => n22910, Z => n22914);
   U11347 : AND2_X1 port map( A1 => n22919, A2 => n22214, ZN => n22578);
   U11348 : AND2_X1 port map( A1 => n22811, A2 => n21199, ZN => n22579);
   U11349 : NOR3_X1 port map( A1 => n22578, A2 => n22579, A3 => n25203, ZN => 
                           n25209);
   U11350 : AND2_X1 port map( A1 => n22919, A2 => n22194, ZN => n22580);
   U11351 : AND2_X1 port map( A1 => n22810, A2 => n21193, ZN => n22581);
   U11352 : NOR3_X1 port map( A1 => n22580, A2 => n22581, A3 => n24499, ZN => 
                           n24505);
   U11353 : AND2_X1 port map( A1 => n22919, A2 => n22209, ZN => n22582);
   U11354 : AND2_X1 port map( A1 => n22803, A2 => n21197, ZN => n22583);
   U11355 : NOR3_X1 port map( A1 => n22582, A2 => n22583, A3 => n25091, ZN => 
                           n25097);
   U11356 : AND2_X1 port map( A1 => n22915, A2 => n22201, ZN => n22584);
   U11357 : AND2_X1 port map( A1 => n22812, A2 => n21188, ZN => n22585);
   U11358 : NOR3_X1 port map( A1 => n22584, A2 => n22585, A3 => n24691, ZN => 
                           n24697);
   U11359 : AND2_X1 port map( A1 => n22911, A2 => n22211, ZN => n22586);
   U11360 : AND2_X1 port map( A1 => n22804, A2 => n21192, ZN => n22587);
   U11361 : NOR3_X1 port map( A1 => n22586, A2 => n22587, A3 => n25155, ZN => 
                           n25161);
   U11362 : AND2_X1 port map( A1 => n22918, A2 => n22219, ZN => n22588);
   U11363 : AND2_X1 port map( A1 => n22809, A2 => n21202, ZN => n22589);
   U11364 : NOR3_X1 port map( A1 => n22588, A2 => n22589, A3 => n25299, ZN => 
                           n25305);
   U11365 : AND2_X1 port map( A1 => n22913, A2 => n22218, ZN => n22590);
   U11366 : AND2_X1 port map( A1 => n22810, A2 => n21180, ZN => n22591);
   U11367 : NOR3_X1 port map( A1 => n22590, A2 => n22591, A3 => n25267, ZN => 
                           n25273);
   U11368 : AND2_X1 port map( A1 => n22917, A2 => n22207, ZN => n22592);
   U11369 : AND2_X1 port map( A1 => n22808, A2 => n21190, ZN => n22593);
   U11370 : NOR3_X1 port map( A1 => n22592, A2 => n22593, A3 => n24851, ZN => 
                           n24857);
   U11371 : AND2_X1 port map( A1 => n22916, A2 => n22217, ZN => n22594);
   U11372 : AND2_X1 port map( A1 => n22808, A2 => n21201, ZN => n22595);
   U11373 : NOR3_X1 port map( A1 => n22594, A2 => n22595, A3 => n25251, ZN => 
                           n25257);
   U11374 : BUF_X1 port map( A => n22910, Z => n22916);
   U11375 : AND2_X1 port map( A1 => n22916, A2 => n22196, ZN => n22596);
   U11376 : AND2_X1 port map( A1 => n22810, A2 => n21185, ZN => n22597);
   U11377 : NOR3_X1 port map( A1 => n22596, A2 => n22597, A3 => n24563, ZN => 
                           n24569);
   U11378 : AND2_X1 port map( A1 => n22914, A2 => n22215, ZN => n22598);
   U11379 : AND2_X1 port map( A1 => n22806, A2 => n21179, ZN => n22599);
   U11380 : NOR3_X1 port map( A1 => n22598, A2 => n22599, A3 => n25219, ZN => 
                           n25225);
   U11381 : AND2_X1 port map( A1 => n22915, A2 => n22193, ZN => n22600);
   U11382 : AND2_X1 port map( A1 => n22808, A2 => n21184, ZN => n22601);
   U11383 : NOR3_X1 port map( A1 => n22600, A2 => n22601, A3 => n24467, ZN => 
                           n24473);
   U11384 : AND2_X1 port map( A1 => n22913, A2 => n22213, ZN => n22602);
   U11385 : AND2_X1 port map( A1 => n22806, A2 => n21198, ZN => n22603);
   U11386 : NOR3_X1 port map( A1 => n22602, A2 => n22603, A3 => n25187, ZN => 
                           n25193);
   U11387 : BUF_X1 port map( A => n22910, Z => n22913);
   U11388 : AND2_X1 port map( A1 => n22915, A2 => n22221, ZN => n22604);
   U11389 : AND2_X1 port map( A1 => n22807, A2 => n21204, ZN => n22605);
   U11390 : NOR3_X1 port map( A1 => n22604, A2 => n22605, A3 => n25331, ZN => 
                           n25337);
   U11391 : BUF_X1 port map( A => n22910, Z => n22915);
   U11392 : AND2_X1 port map( A1 => n22911, A2 => n22192, ZN => n22606);
   U11393 : AND2_X1 port map( A1 => n22812, A2 => n21174, ZN => n22607);
   U11394 : NOR3_X1 port map( A1 => n22606, A2 => n22607, A3 => n24451, ZN => 
                           n24457);
   U11395 : BUF_X1 port map( A => n22910, Z => n22911);
   U11396 : AND2_X1 port map( A1 => n22915, A2 => n22205, ZN => n22608);
   U11397 : AND2_X1 port map( A1 => n22805, A2 => n21196, ZN => n22609);
   U11398 : NOR3_X1 port map( A1 => n22608, A2 => n22609, A3 => n24819, ZN => 
                           n24825);
   U11399 : AND2_X1 port map( A1 => n22912, A2 => n22212, ZN => n22610);
   U11400 : AND2_X1 port map( A1 => n22810, A2 => n21178, ZN => n22611);
   U11401 : NOR3_X1 port map( A1 => n22610, A2 => n22611, A3 => n25171, ZN => 
                           n25177);
   U11402 : AND2_X1 port map( A1 => n22916, A2 => n22220, ZN => n22612);
   U11403 : AND2_X1 port map( A1 => n22808, A2 => n21181, ZN => n22613);
   U11404 : NOR3_X1 port map( A1 => n22612, A2 => n22613, A3 => n25315, ZN => 
                           n25321);
   U11405 : AND2_X1 port map( A1 => n22911, A2 => n22190, ZN => n22614);
   U11406 : AND2_X1 port map( A1 => n22807, A2 => n21182, ZN => n22615);
   U11407 : NOR3_X1 port map( A1 => n22614, A2 => n22615, A3 => n24403, ZN => 
                           n24409);
   U11408 : AND2_X1 port map( A1 => n22910, A2 => n22195, ZN => n22616);
   U11409 : AND2_X1 port map( A1 => n22803, A2 => n21207, ZN => n22617);
   U11410 : NOR3_X1 port map( A1 => n22616, A2 => n22617, A3 => n24515, ZN => 
                           n24521);
   U11411 : AND2_X1 port map( A1 => n22913, A2 => n22197, ZN => n22618);
   U11412 : AND2_X1 port map( A1 => n22809, A2 => n21194, ZN => n22619);
   U11413 : NOR3_X1 port map( A1 => n22618, A2 => n22619, A3 => n24579, ZN => 
                           n24585);
   U11414 : AND2_X1 port map( A1 => n22913, A2 => n22206, ZN => n22620);
   U11415 : AND2_X1 port map( A1 => n22806, A2 => n21189, ZN => n22621);
   U11416 : NOR3_X1 port map( A1 => n22620, A2 => n22621, A3 => n24835, ZN => 
                           n24841);
   U11417 : AND2_X1 port map( A1 => n22915, A2 => n22216, ZN => n22622);
   U11418 : AND2_X1 port map( A1 => n22812, A2 => n21200, ZN => n22623);
   U11419 : NOR3_X1 port map( A1 => n22622, A2 => n22623, A3 => n25235, ZN => 
                           n25241);
   U11420 : AND2_X1 port map( A1 => n22917, A2 => n22208, ZN => n22624);
   U11421 : AND2_X1 port map( A1 => n22807, A2 => n21191, ZN => n22625);
   U11422 : NOR3_X1 port map( A1 => n22624, A2 => n22625, A3 => n24979, ZN => 
                           n24985);
   U11423 : NAND3_X1 port map( A1 => n24087, A2 => n22512, A3 => n21415, ZN => 
                           n22628);
   U11424 : AND2_X1 port map( A1 => n22911, A2 => n22200, ZN => n22626);
   U11425 : AND2_X1 port map( A1 => n22809, A2 => n21187, ZN => n22627);
   U11426 : NOR3_X1 port map( A1 => n22626, A2 => n22627, A3 => n24627, ZN => 
                           n24633);
   U11427 : BUF_X1 port map( A => n22930, Z => n22640);
   U11428 : BUF_X1 port map( A => n22931, Z => n22643);
   U11429 : BUF_X1 port map( A => n22675, Z => n22646);
   U11430 : BUF_X1 port map( A => n22949, Z => n22649);
   U11431 : CLKBUF_X1 port map( A => n22948, Z => n22629);
   U11432 : BUF_X1 port map( A => n22948, Z => n22630);
   U11433 : BUF_X1 port map( A => n22948, Z => n22631);
   U11434 : CLKBUF_X1 port map( A => n22950, Z => n22632);
   U11435 : BUF_X1 port map( A => n22950, Z => n22633);
   U11436 : BUF_X1 port map( A => n22950, Z => n22634);
   U11437 : CLKBUF_X3 port map( A => n25387, Z => n22635);
   U11438 : CLKBUF_X3 port map( A => n25387, Z => n22636);
   U11439 : CLKBUF_X3 port map( A => n25387, Z => n22637);
   U11440 : CLKBUF_X3 port map( A => n25387, Z => n22638);
   U11441 : BUF_X1 port map( A => n22930, Z => n22641);
   U11442 : BUF_X1 port map( A => n22930, Z => n22642);
   U11443 : BUF_X1 port map( A => n22931, Z => n22644);
   U11444 : BUF_X1 port map( A => n22931, Z => n22645);
   U11445 : BUF_X1 port map( A => n22675, Z => n22647);
   U11446 : BUF_X1 port map( A => n22675, Z => n22648);
   U11447 : BUF_X1 port map( A => n22949, Z => n22650);
   U11448 : BUF_X1 port map( A => n22949, Z => n22651);
   U11449 : AOI22_X2 port map( A1 => MEM_BUSread(55), A2 => n23052, B1 => 
                           DATAIN(55), B2 => n23040, ZN => n16605);
   U11450 : AOI22_X2 port map( A1 => MEM_BUSread(31), A2 => n23051, B1 => 
                           DATAIN(31), B2 => n23041, ZN => n16617);
   U11451 : AOI22_X2 port map( A1 => MEM_BUSread(5), A2 => n23050, B1 => 
                           DATAIN(5), B2 => n23042, ZN => n16630);
   U11452 : AOI22_X2 port map( A1 => MEM_BUSread(14), A2 => n23049, B1 => 
                           DATAIN(14), B2 => n23043, ZN => n16640);
   U11453 : AOI22_X2 port map( A1 => MEM_BUSread(38), A2 => n23048, B1 => 
                           DATAIN(38), B2 => n23044, ZN => n16652);
   U11454 : AOI22_X2 port map( A1 => MEM_BUSread(53), A2 => n23052, B1 => 
                           DATAIN(53), B2 => n23040, ZN => n16606);
   U11455 : AOI22_X2 port map( A1 => MEM_BUSread(29), A2 => n23051, B1 => 
                           DATAIN(29), B2 => n23041, ZN => n16618);
   U11456 : AOI22_X2 port map( A1 => MEM_BUSread(3), A2 => n23050, B1 => 
                           DATAIN(3), B2 => n23042, ZN => n16631);
   U11457 : AOI22_X2 port map( A1 => MEM_BUSread(16), A2 => n23049, B1 => 
                           DATAIN(16), B2 => n23043, ZN => n16641);
   U11458 : AOI22_X2 port map( A1 => MEM_BUSread(40), A2 => n23048, B1 => 
                           DATAIN(40), B2 => n23044, ZN => n16653);
   U11459 : AOI22_X2 port map( A1 => MEM_BUSread(51), A2 => n23052, B1 => 
                           DATAIN(51), B2 => n23040, ZN => n16607);
   U11460 : AOI22_X2 port map( A1 => MEM_BUSread(27), A2 => n23051, B1 => 
                           DATAIN(27), B2 => n23041, ZN => n16619);
   U11461 : AOI22_X2 port map( A1 => MEM_BUSread(1), A2 => n23050, B1 => 
                           DATAIN(1), B2 => n23042, ZN => n16632);
   U11462 : AOI22_X2 port map( A1 => MEM_BUSread(18), A2 => n23049, B1 => 
                           DATAIN(18), B2 => n23043, ZN => n16642);
   U11463 : AOI22_X2 port map( A1 => MEM_BUSread(42), A2 => n23048, B1 => 
                           DATAIN(42), B2 => n23044, ZN => n16654);
   U11464 : AOI22_X2 port map( A1 => MEM_BUSread(49), A2 => n23052, B1 => 
                           DATAIN(49), B2 => n23040, ZN => n16608);
   U11465 : AOI22_X2 port map( A1 => MEM_BUSread(25), A2 => n23051, B1 => 
                           DATAIN(25), B2 => n23041, ZN => n16620);
   U11466 : AOI22_X2 port map( A1 => MEM_BUSread(2), A2 => n23050, B1 => 
                           DATAIN(2), B2 => n23042, ZN => n16634);
   U11467 : AOI22_X2 port map( A1 => MEM_BUSread(20), A2 => n23049, B1 => 
                           DATAIN(20), B2 => n23043, ZN => n16643);
   U11468 : AOI22_X2 port map( A1 => MEM_BUSread(44), A2 => n23048, B1 => 
                           DATAIN(44), B2 => n23044, ZN => n16655);
   U11469 : AOI22_X2 port map( A1 => MEM_BUSread(47), A2 => n23052, B1 => 
                           DATAIN(47), B2 => n23040, ZN => n16609);
   U11470 : AOI22_X2 port map( A1 => MEM_BUSread(23), A2 => n23051, B1 => 
                           DATAIN(23), B2 => n23041, ZN => n16621);
   U11471 : AOI22_X2 port map( A1 => MEM_BUSread(4), A2 => n23050, B1 => 
                           DATAIN(4), B2 => n23042, ZN => n16635);
   U11472 : AOI22_X2 port map( A1 => MEM_BUSread(22), A2 => n23049, B1 => 
                           DATAIN(22), B2 => n23043, ZN => n16644);
   U11473 : AOI22_X2 port map( A1 => MEM_BUSread(46), A2 => n23048, B1 => 
                           DATAIN(46), B2 => n23044, ZN => n16656);
   U11474 : AOI22_X2 port map( A1 => MEM_BUSread(45), A2 => n23052, B1 => 
                           DATAIN(45), B2 => n23040, ZN => n16610);
   U11475 : AOI22_X2 port map( A1 => MEM_BUSread(21), A2 => n23051, B1 => 
                           DATAIN(21), B2 => n23041, ZN => n16622);
   U11476 : AOI22_X2 port map( A1 => MEM_BUSread(24), A2 => n23049, B1 => 
                           DATAIN(24), B2 => n23043, ZN => n16645);
   U11477 : AOI22_X2 port map( A1 => MEM_BUSread(48), A2 => n23048, B1 => 
                           DATAIN(48), B2 => n23044, ZN => n16657);
   U11478 : AOI22_X2 port map( A1 => MEM_BUSread(7), A2 => n23050, B1 => 
                           DATAIN(7), B2 => n23042, ZN => n16629);
   U11479 : AOI22_X2 port map( A1 => MEM_BUSread(43), A2 => n23052, B1 => 
                           DATAIN(43), B2 => n23040, ZN => n16611);
   U11480 : AOI22_X2 port map( A1 => MEM_BUSread(19), A2 => n23051, B1 => 
                           DATAIN(19), B2 => n23041, ZN => n16623);
   U11481 : AOI22_X2 port map( A1 => MEM_BUSread(26), A2 => n23049, B1 => 
                           DATAIN(26), B2 => n23043, ZN => n16646);
   U11482 : AOI22_X2 port map( A1 => MEM_BUSread(50), A2 => n23048, B1 => 
                           DATAIN(50), B2 => n23044, ZN => n16658);
   U11483 : AOI22_X2 port map( A1 => MEM_BUSread(0), A2 => n23050, B1 => 
                           DATAIN(0), B2 => n23042, ZN => n16633);
   U11484 : CLKBUF_X3 port map( A => n25381, Z => n22652);
   U11485 : NAND2_X2 port map( A1 => n22698, A2 => n22699, ZN => n25381);
   U11486 : BUF_X2 port map( A => n25392, Z => n22947);
   U11487 : INV_X2 port map( A => n23032, ZN => n23031);
   U11488 : BUF_X1 port map( A => n23520, Z => n23517);
   U11489 : BUF_X1 port map( A => n23520, Z => n23518);
   U11490 : BUF_X1 port map( A => n23520, Z => n23519);
   U11491 : BUF_X1 port map( A => n23529, Z => n23527);
   U11492 : BUF_X1 port map( A => n23549, Z => n23547);
   U11493 : BUF_X1 port map( A => n23569, Z => n23567);
   U11494 : BUF_X1 port map( A => n23589, Z => n23587);
   U11495 : BUF_X1 port map( A => n23539, Z => n23537);
   U11496 : BUF_X1 port map( A => n23579, Z => n23577);
   U11497 : BUF_X1 port map( A => n23559, Z => n23557);
   U11498 : BUF_X1 port map( A => n23529, Z => n23528);
   U11499 : BUF_X1 port map( A => n23549, Z => n23548);
   U11500 : BUF_X1 port map( A => n23569, Z => n23568);
   U11501 : BUF_X1 port map( A => n23589, Z => n23588);
   U11502 : BUF_X1 port map( A => n23539, Z => n23538);
   U11503 : BUF_X1 port map( A => n23579, Z => n23578);
   U11504 : BUF_X1 port map( A => n23559, Z => n23558);
   U11505 : BUF_X1 port map( A => n23609, Z => n23607);
   U11506 : BUF_X1 port map( A => n23629, Z => n23627);
   U11507 : BUF_X1 port map( A => n23649, Z => n23647);
   U11508 : BUF_X1 port map( A => n23669, Z => n23667);
   U11509 : BUF_X1 port map( A => n23609, Z => n23608);
   U11510 : BUF_X1 port map( A => n23629, Z => n23628);
   U11511 : BUF_X1 port map( A => n23649, Z => n23648);
   U11512 : BUF_X1 port map( A => n23669, Z => n23668);
   U11513 : BUF_X1 port map( A => n23659, Z => n23657);
   U11514 : BUF_X1 port map( A => n23659, Z => n23658);
   U11515 : BUF_X1 port map( A => n23599, Z => n23597);
   U11516 : BUF_X1 port map( A => n23619, Z => n23617);
   U11517 : BUF_X1 port map( A => n23639, Z => n23637);
   U11518 : BUF_X1 port map( A => n23599, Z => n23598);
   U11519 : BUF_X1 port map( A => n23619, Z => n23618);
   U11520 : BUF_X1 port map( A => n23639, Z => n23638);
   U11521 : BUF_X1 port map( A => n23529, Z => n23526);
   U11522 : BUF_X1 port map( A => n23549, Z => n23546);
   U11523 : BUF_X1 port map( A => n23569, Z => n23566);
   U11524 : BUF_X1 port map( A => n23589, Z => n23586);
   U11525 : BUF_X1 port map( A => n23539, Z => n23536);
   U11526 : BUF_X1 port map( A => n23559, Z => n23556);
   U11527 : BUF_X1 port map( A => n23579, Z => n23576);
   U11528 : BUF_X1 port map( A => n23609, Z => n23606);
   U11529 : BUF_X1 port map( A => n23629, Z => n23626);
   U11530 : BUF_X1 port map( A => n23649, Z => n23646);
   U11531 : BUF_X1 port map( A => n23669, Z => n23666);
   U11532 : BUF_X1 port map( A => n23659, Z => n23656);
   U11533 : BUF_X1 port map( A => n23599, Z => n23596);
   U11534 : BUF_X1 port map( A => n23619, Z => n23616);
   U11535 : BUF_X1 port map( A => n23639, Z => n23636);
   U11536 : BUF_X1 port map( A => n22653, Z => n23355);
   U11537 : BUF_X1 port map( A => n22653, Z => n23354);
   U11538 : BUF_X1 port map( A => n23330, Z => n23329);
   U11539 : BUF_X1 port map( A => n22654, Z => n23371);
   U11540 : BUF_X1 port map( A => n22654, Z => n23370);
   U11541 : BUF_X1 port map( A => n22655, Z => n23363);
   U11542 : BUF_X1 port map( A => n22655, Z => n23362);
   U11543 : BUF_X1 port map( A => n23330, Z => n23328);
   U11544 : BUF_X1 port map( A => n23319, Z => n23317);
   U11545 : BUF_X1 port map( A => n23319, Z => n23316);
   U11546 : BUF_X1 port map( A => n23319, Z => n23318);
   U11547 : BUF_X1 port map( A => n23307, Z => n23305);
   U11548 : BUF_X1 port map( A => n23307, Z => n23306);
   U11549 : BUF_X1 port map( A => n23296, Z => n23294);
   U11550 : BUF_X1 port map( A => n23296, Z => n23293);
   U11551 : BUF_X1 port map( A => n23296, Z => n23295);
   U11552 : BUF_X1 port map( A => n22656, Z => n23388);
   U11553 : BUF_X1 port map( A => n22656, Z => n23387);
   U11554 : BUF_X1 port map( A => n22657, Z => n23396);
   U11555 : BUF_X1 port map( A => n22657, Z => n23395);
   U11556 : BUF_X1 port map( A => n22658, Z => n23404);
   U11557 : BUF_X1 port map( A => n22658, Z => n23403);
   U11558 : BUF_X1 port map( A => n22659, Z => n23339);
   U11559 : BUF_X1 port map( A => n22659, Z => n23338);
   U11560 : BUF_X1 port map( A => n22660, Z => n23267);
   U11561 : BUF_X1 port map( A => n22660, Z => n23266);
   U11562 : BUF_X1 port map( A => n23372, Z => n23380);
   U11563 : BUF_X1 port map( A => n23372, Z => n23379);
   U11564 : BUF_X1 port map( A => n22661, Z => n23347);
   U11565 : BUF_X1 port map( A => n22661, Z => n23346);
   U11566 : BUF_X1 port map( A => n22662, Z => n23259);
   U11567 : BUF_X1 port map( A => n22662, Z => n23258);
   U11568 : BUF_X1 port map( A => n22663, Z => n23251);
   U11569 : BUF_X1 port map( A => n22663, Z => n23250);
   U11570 : BUF_X1 port map( A => n21448, Z => n23227);
   U11571 : BUF_X1 port map( A => n21448, Z => n23226);
   U11572 : BUF_X1 port map( A => n21450, Z => n23235);
   U11573 : BUF_X1 port map( A => n21450, Z => n23234);
   U11574 : BUF_X1 port map( A => n21451, Z => n23219);
   U11575 : BUF_X1 port map( A => n21451, Z => n23218);
   U11576 : BUF_X1 port map( A => n21452, Z => n23243);
   U11577 : BUF_X1 port map( A => n21452, Z => n23242);
   U11578 : BUF_X1 port map( A => n23425, Z => n23424);
   U11579 : BUF_X1 port map( A => n23469, Z => n23468);
   U11580 : BUF_X1 port map( A => n23480, Z => n23479);
   U11581 : BUF_X1 port map( A => n23512, Z => n23510);
   U11582 : BUF_X1 port map( A => n23512, Z => n23509);
   U11583 : BUF_X1 port map( A => n23414, Z => n23413);
   U11584 : BUF_X1 port map( A => n23414, Z => n23412);
   U11585 : BUF_X1 port map( A => n23469, Z => n23467);
   U11586 : BUF_X1 port map( A => n23469, Z => n23466);
   U11587 : BUF_X1 port map( A => n23425, Z => n23423);
   U11588 : BUF_X1 port map( A => n23480, Z => n23478);
   U11589 : BUF_X1 port map( A => n23480, Z => n23477);
   U11590 : BUF_X1 port map( A => n23457, Z => n23455);
   U11591 : BUF_X1 port map( A => n23457, Z => n23454);
   U11592 : BUF_X1 port map( A => n23496, Z => n23494);
   U11593 : BUF_X1 port map( A => n23496, Z => n23493);
   U11594 : BUF_X1 port map( A => n23441, Z => n23439);
   U11595 : BUF_X1 port map( A => n23441, Z => n23438);
   U11596 : BUF_X1 port map( A => n22677, Z => n22992);
   U11597 : AND2_X1 port map( A1 => n23027, A2 => n23036, ZN => n22676);
   U11598 : BUF_X1 port map( A => n24285, Z => n23183);
   U11599 : BUF_X1 port map( A => n24285, Z => n23182);
   U11600 : BUF_X1 port map( A => n24281, Z => n23151);
   U11601 : BUF_X1 port map( A => n24281, Z => n23150);
   U11602 : BUF_X1 port map( A => n23521, Z => n23520);
   U11603 : BUF_X1 port map( A => n24142, Z => n23086);
   U11604 : BUF_X1 port map( A => n24142, Z => n23087);
   U11605 : BUF_X1 port map( A => n24277, Z => n23119);
   U11606 : BUF_X1 port map( A => n24277, Z => n23118);
   U11607 : BUF_X1 port map( A => n24140, Z => n23078);
   U11608 : BUF_X1 port map( A => n24140, Z => n23079);
   U11609 : BUF_X1 port map( A => n24276, Z => n23111);
   U11610 : BUF_X1 port map( A => n24276, Z => n23110);
   U11611 : BUF_X1 port map( A => n24274, Z => n23095);
   U11612 : BUF_X1 port map( A => n24274, Z => n23094);
   U11613 : BUF_X1 port map( A => n24278, Z => n23127);
   U11614 : BUF_X1 port map( A => n24278, Z => n23126);
   U11615 : BUF_X1 port map( A => n24275, Z => n23103);
   U11616 : BUF_X1 port map( A => n24275, Z => n23102);
   U11617 : BUF_X1 port map( A => n24279, Z => n23135);
   U11618 : BUF_X1 port map( A => n24279, Z => n23134);
   U11619 : BUF_X1 port map( A => n24283, Z => n23167);
   U11620 : BUF_X1 port map( A => n24283, Z => n23166);
   U11621 : BUF_X1 port map( A => n23531, Z => n23529);
   U11622 : BUF_X1 port map( A => n23551, Z => n23549);
   U11623 : BUF_X1 port map( A => n23571, Z => n23569);
   U11624 : BUF_X1 port map( A => n23591, Z => n23589);
   U11625 : BUF_X1 port map( A => n23541, Z => n23539);
   U11626 : BUF_X1 port map( A => n23581, Z => n23579);
   U11627 : BUF_X1 port map( A => n23561, Z => n23559);
   U11628 : BUF_X1 port map( A => n24280, Z => n23143);
   U11629 : BUF_X1 port map( A => n24280, Z => n23142);
   U11630 : BUF_X1 port map( A => n24137, Z => n23070);
   U11631 : BUF_X1 port map( A => n24137, Z => n23071);
   U11632 : BUF_X1 port map( A => n23748, Z => n23756);
   U11633 : BUF_X1 port map( A => n23748, Z => n23755);
   U11634 : BUF_X1 port map( A => n23611, Z => n23609);
   U11635 : BUF_X1 port map( A => n23631, Z => n23629);
   U11636 : BUF_X1 port map( A => n23651, Z => n23649);
   U11637 : BUF_X1 port map( A => n23671, Z => n23669);
   U11638 : BUF_X1 port map( A => n23661, Z => n23659);
   U11639 : BUF_X1 port map( A => n23601, Z => n23599);
   U11640 : BUF_X1 port map( A => n23621, Z => n23619);
   U11641 : BUF_X1 port map( A => n23641, Z => n23639);
   U11642 : BUF_X1 port map( A => n23590, Z => n23585);
   U11643 : BUF_X1 port map( A => n23550, Z => n23545);
   U11644 : BUF_X1 port map( A => n23530, Z => n23525);
   U11645 : BUF_X1 port map( A => n23570, Z => n23565);
   U11646 : BUF_X1 port map( A => n23540, Z => n23535);
   U11647 : BUF_X1 port map( A => n23560, Z => n23555);
   U11648 : BUF_X1 port map( A => n23580, Z => n23575);
   U11649 : BUF_X1 port map( A => n23650, Z => n23645);
   U11650 : BUF_X1 port map( A => n23670, Z => n23665);
   U11651 : BUF_X1 port map( A => n23610, Z => n23605);
   U11652 : BUF_X1 port map( A => n23630, Z => n23625);
   U11653 : BUF_X1 port map( A => n23660, Z => n23655);
   U11654 : BUF_X1 port map( A => n23722, Z => n23730);
   U11655 : BUF_X1 port map( A => n23722, Z => n23729);
   U11656 : BUF_X1 port map( A => n15212, Z => n23764);
   U11657 : BUF_X1 port map( A => n15212, Z => n23763);
   U11658 : BUF_X1 port map( A => n23640, Z => n23635);
   U11659 : BUF_X1 port map( A => n23600, Z => n23595);
   U11660 : BUF_X1 port map( A => n23620, Z => n23615);
   U11661 : BUF_X1 port map( A => n15211, Z => n23772);
   U11662 : BUF_X1 port map( A => n15211, Z => n23771);
   U11663 : BUF_X1 port map( A => n23790, Z => n23798);
   U11664 : BUF_X1 port map( A => n23790, Z => n23797);
   U11665 : BUF_X1 port map( A => n23713, Z => n23721);
   U11666 : BUF_X1 port map( A => n23713, Z => n23720);
   U11667 : BUF_X1 port map( A => n22664, Z => n23806);
   U11668 : BUF_X1 port map( A => n22664, Z => n23805);
   U11669 : BUF_X1 port map( A => n23781, Z => n23789);
   U11670 : BUF_X1 port map( A => n23781, Z => n23788);
   U11671 : BUF_X1 port map( A => n23696, Z => n23704);
   U11672 : BUF_X1 port map( A => n23696, Z => n23703);
   U11673 : BUF_X1 port map( A => n22665, Z => n23780);
   U11674 : BUF_X1 port map( A => n22665, Z => n23779);
   U11675 : BUF_X1 port map( A => n22666, Z => n23712);
   U11676 : BUF_X1 port map( A => n22666, Z => n23711);
   U11677 : AND2_X1 port map( A1 => n21445, A2 => n23424, ZN => n22653);
   U11678 : BUF_X1 port map( A => n23739, Z => n23747);
   U11679 : BUF_X1 port map( A => n23739, Z => n23746);
   U11680 : BUF_X1 port map( A => n22682, Z => n23330);
   U11681 : AND2_X1 port map( A1 => n21445, A2 => n23479, ZN => n22654);
   U11682 : AND2_X1 port map( A1 => n21445, A2 => n23468, ZN => n22655);
   U11683 : BUF_X1 port map( A => n15221, Z => n23695);
   U11684 : BUF_X1 port map( A => n15221, Z => n23694);
   U11685 : BUF_X1 port map( A => n22683, Z => n23319);
   U11686 : BUF_X1 port map( A => n22680, Z => n23307);
   U11687 : BUF_X1 port map( A => n22679, Z => n23296);
   U11688 : BUF_X1 port map( A => n23847, Z => n23845);
   U11689 : BUF_X1 port map( A => n23847, Z => n23844);
   U11690 : BUF_X1 port map( A => n23331, Z => n23327);
   U11691 : BUF_X1 port map( A => n23320, Z => n23315);
   U11692 : BUF_X1 port map( A => n23308, Z => n23304);
   U11693 : BUF_X1 port map( A => n23297, Z => n23292);
   U11694 : NAND2_X1 port map( A1 => n21445, A2 => n23443, ZN => n22656);
   U11695 : NAND2_X1 port map( A1 => n21445, A2 => n23427, ZN => n22657);
   U11696 : NAND2_X1 port map( A1 => n21445, A2 => n23482, ZN => n22658);
   U11697 : BUF_X1 port map( A => n23831, Z => n23828);
   U11698 : BUF_X1 port map( A => n23831, Z => n23829);
   U11699 : BUF_X1 port map( A => n15215, Z => n23738);
   U11700 : BUF_X1 port map( A => n15215, Z => n23737);
   U11701 : BUF_X1 port map( A => n23879, Z => n23877);
   U11702 : BUF_X1 port map( A => n23879, Z => n23876);
   U11703 : NAND2_X1 port map( A1 => n23491, A2 => n21447, ZN => n22659);
   U11704 : NAND2_X1 port map( A1 => n23452, A2 => n21447, ZN => n22660);
   U11705 : BUF_X1 port map( A => n16795, Z => n23372);
   U11706 : NAND2_X1 port map( A1 => n21445, A2 => n23413, ZN => n22661);
   U11707 : BUF_X1 port map( A => n15223, Z => n23679);
   U11708 : BUF_X1 port map( A => n15223, Z => n23678);
   U11709 : BUF_X1 port map( A => n15222, Z => n23687);
   U11710 : BUF_X1 port map( A => n15222, Z => n23686);
   U11711 : NAND2_X1 port map( A1 => n21447, A2 => n23424, ZN => n22662);
   U11712 : NAND2_X1 port map( A1 => n21447, A2 => n23479, ZN => n22663);
   U11713 : BUF_X1 port map( A => n23863, Z => n23861);
   U11714 : BUF_X1 port map( A => n23863, Z => n23860);
   U11715 : BUF_X1 port map( A => n22667, Z => n23512);
   U11716 : BUF_X1 port map( A => n22668, Z => n23457);
   U11717 : BUF_X1 port map( A => n22669, Z => n23441);
   U11718 : BUF_X1 port map( A => n22670, Z => n23496);
   U11719 : BUF_X1 port map( A => n23458, Z => n23453);
   U11720 : BUF_X1 port map( A => n23497, Z => n23492);
   U11721 : BUF_X1 port map( A => n23513, Z => n23508);
   U11722 : BUF_X1 port map( A => n22684, Z => n23425);
   U11723 : BUF_X1 port map( A => n23442, Z => n23437);
   U11724 : BUF_X1 port map( A => n22685, Z => n23469);
   U11725 : BUF_X1 port map( A => n22686, Z => n23480);
   U11726 : BUF_X1 port map( A => n22687, Z => n23414);
   U11727 : BUF_X1 port map( A => n23415, Z => n23411);
   U11728 : BUF_X1 port map( A => n23470, Z => n23465);
   U11729 : BUF_X1 port map( A => n23426, Z => n23422);
   U11730 : BUF_X1 port map( A => n23481, Z => n23476);
   U11731 : AND2_X1 port map( A1 => n23984, A2 => n23983, ZN => n22677);
   U11732 : BUF_X1 port map( A => n22681, Z => n22998);
   U11733 : BUF_X1 port map( A => n24282, Z => n23159);
   U11734 : BUF_X1 port map( A => n24282, Z => n23158);
   U11735 : BUF_X1 port map( A => n24284, Z => n23175);
   U11736 : BUF_X1 port map( A => n24284, Z => n23174);
   U11737 : BUF_X1 port map( A => n16725, Z => n23591);
   U11738 : BUF_X1 port map( A => n16734, Z => n23531);
   U11739 : BUF_X1 port map( A => n16732, Z => n23551);
   U11740 : BUF_X1 port map( A => n16730, Z => n23571);
   U11741 : BUF_X1 port map( A => n16733, Z => n23541);
   U11742 : BUF_X1 port map( A => n16731, Z => n23561);
   U11743 : BUF_X1 port map( A => n16728, Z => n23581);
   U11744 : BUF_X1 port map( A => n23832, Z => n23827);
   U11745 : BUF_X1 port map( A => n15213, Z => n23748);
   U11746 : BUF_X1 port map( A => n16718, Z => n23651);
   U11747 : BUF_X1 port map( A => n16713, Z => n23671);
   U11748 : BUF_X1 port map( A => n16722, Z => n23611);
   U11749 : BUF_X1 port map( A => n16720, Z => n23631);
   U11750 : BUF_X1 port map( A => n16716, Z => n23661);
   U11751 : BUF_X1 port map( A => n16719, Z => n23641);
   U11752 : BUF_X1 port map( A => n16724, Z => n23601);
   U11753 : BUF_X1 port map( A => n16721, Z => n23621);
   U11754 : BUF_X1 port map( A => n21440, Z => n23847);
   U11755 : BUF_X1 port map( A => n15217, Z => n23722);
   U11756 : BUF_X1 port map( A => n15207, Z => n23790);
   U11757 : BUF_X1 port map( A => n15218, Z => n23713);
   U11758 : NAND2_X1 port map( A1 => n16552, A2 => n23849, ZN => n22664);
   U11759 : BUF_X1 port map( A => n15208, Z => n23781);
   U11760 : BUF_X1 port map( A => n23848, Z => n23843);
   U11761 : BUF_X1 port map( A => n15220, Z => n23696);
   U11762 : NAND2_X1 port map( A1 => n16552, A2 => n23865, ZN => n22665);
   U11763 : BUF_X1 port map( A => n23864, Z => n23859);
   U11764 : BUF_X1 port map( A => n21443, Z => n23863);
   U11765 : BUF_X1 port map( A => n21444, Z => n23879);
   U11766 : AND2_X1 port map( A1 => n23826, A2 => n16555, ZN => n22666);
   U11767 : BUF_X1 port map( A => n15214, Z => n23739);
   U11768 : BUF_X1 port map( A => n23880, Z => n23875);
   U11769 : BUF_X1 port map( A => n21438, Z => n23831);
   U11770 : BUF_X1 port map( A => n23881, Z => n23889);
   U11771 : BUF_X1 port map( A => n23881, Z => n23888);
   U11772 : BUF_X1 port map( A => n23807, Z => n23815);
   U11773 : BUF_X1 port map( A => n23807, Z => n23814);
   U11774 : NOR3_X1 port map( A1 => n18526, A2 => n25401, A3 => n25402, ZN => 
                           n22667);
   U11775 : NOR3_X1 port map( A1 => n18525, A2 => n18526, A3 => n25402, ZN => 
                           n22668);
   U11776 : NOR3_X1 port map( A1 => n18525, A2 => n25400, A3 => n25402, ZN => 
                           n22669);
   U11777 : NOR3_X1 port map( A1 => n25400, A2 => n25401, A3 => n25402, ZN => 
                           n22670);
   U11778 : BUF_X1 port map( A => n23195, Z => n23203);
   U11779 : BUF_X1 port map( A => n23195, Z => n23202);
   U11780 : BUF_X1 port map( A => n21454, Z => n23211);
   U11781 : BUF_X1 port map( A => n21454, Z => n23210);
   U11782 : AND2_X1 port map( A1 => n22990, A2 => n20834, ZN => n22681);
   U11783 : BUF_X1 port map( A => n23934, Z => n23933);
   U11784 : BUF_X1 port map( A => n23934, Z => n23932);
   U11785 : BUF_X1 port map( A => n23272, Z => n23271);
   U11786 : BUF_X1 port map( A => n21459, Z => n23193);
   U11787 : BUF_X1 port map( A => n21459, Z => n23194);
   U11788 : CLKBUF_X3 port map( A => n25381, Z => n22933);
   U11789 : BUF_X1 port map( A => n24135, Z => n23062);
   U11790 : BUF_X1 port map( A => n24135, Z => n23063);
   U11791 : XNOR2_X1 port map( A => n22692, B => n24159, ZN => n25402);
   U11792 : NAND2_X1 port map( A1 => n23992, A2 => n22529, ZN => n22671);
   U11793 : BUF_X1 port map( A => n23273, Z => n23272);
   U11794 : BUF_X1 port map( A => n21457, Z => n23054);
   U11795 : BUF_X1 port map( A => n23908, Z => n23916);
   U11796 : BUF_X1 port map( A => n23908, Z => n23915);
   U11797 : BUF_X1 port map( A => n23917, Z => n23925);
   U11798 : BUF_X1 port map( A => n23917, Z => n23924);
   U11799 : BUF_X1 port map( A => n22672, Z => n23942);
   U11800 : BUF_X1 port map( A => n22672, Z => n23941);
   U11801 : BUF_X1 port map( A => n23907, Z => n23906);
   U11802 : BUF_X1 port map( A => n23907, Z => n23905);
   U11803 : BUF_X1 port map( A => n21458, Z => n23046);
   U11804 : BUF_X1 port map( A => n21458, Z => n23047);
   U11805 : BUF_X1 port map( A => n21457, Z => n23055);
   U11806 : BUF_X1 port map( A => n23898, Z => n23897);
   U11807 : BUF_X1 port map( A => n23898, Z => n23896);
   U11808 : BUF_X1 port map( A => n24095, Z => n23022);
   U11809 : BUF_X1 port map( A => n22766, Z => n23946);
   U11810 : BUF_X1 port map( A => n22767, Z => n23005);
   U11811 : BUF_X1 port map( A => n24127, Z => n23038);
   U11812 : AND2_X1 port map( A1 => n25407, A2 => ADD_RD2(2), ZN => n22672);
   U11813 : INV_X1 port map( A => n22673, ZN => n22674);
   U11814 : BUF_X1 port map( A => n25384, Z => n22675);
   U11815 : INV_X1 port map( A => n23517, ZN => n23515);
   U11816 : INV_X1 port map( A => n23517, ZN => n23514);
   U11817 : BUF_X1 port map( A => n23518, Z => n22813);
   U11818 : BUF_X1 port map( A => n23518, Z => n22814);
   U11819 : BUF_X1 port map( A => n23518, Z => n22815);
   U11820 : BUF_X1 port map( A => n23519, Z => n22816);
   U11821 : BUF_X1 port map( A => n23519, Z => n22817);
   U11822 : BUF_X1 port map( A => n23519, Z => n22818);
   U11823 : INV_X1 port map( A => n22992, ZN => n22990);
   U11824 : INV_X1 port map( A => n23526, ZN => n23522);
   U11825 : INV_X1 port map( A => n23546, ZN => n23542);
   U11826 : INV_X1 port map( A => n23566, ZN => n23562);
   U11827 : INV_X1 port map( A => n23586, ZN => n23582);
   U11828 : INV_X1 port map( A => n23536, ZN => n23532);
   U11829 : INV_X1 port map( A => n23556, ZN => n23552);
   U11830 : INV_X1 port map( A => n23576, ZN => n23572);
   U11831 : INV_X1 port map( A => n23306, ZN => n23298);
   U11832 : INV_X1 port map( A => n23329, ZN => n23321);
   U11833 : INV_X1 port map( A => n23329, ZN => n23322);
   U11834 : INV_X1 port map( A => n23306, ZN => n23299);
   U11835 : INV_X1 port map( A => n23295, ZN => n23286);
   U11836 : INV_X1 port map( A => n23318, ZN => n23309);
   U11837 : INV_X1 port map( A => n23318, ZN => n23310);
   U11838 : INV_X1 port map( A => n23295, ZN => n23287);
   U11839 : INV_X1 port map( A => n23606, ZN => n23602);
   U11840 : INV_X1 port map( A => n23626, ZN => n23622);
   U11841 : INV_X1 port map( A => n23646, ZN => n23642);
   U11842 : INV_X1 port map( A => n23666, ZN => n23662);
   U11843 : INV_X1 port map( A => n23328, ZN => n23323);
   U11844 : INV_X1 port map( A => n23328, ZN => n23324);
   U11845 : INV_X1 port map( A => n23305, ZN => n23300);
   U11846 : INV_X1 port map( A => n23305, ZN => n23301);
   U11847 : INV_X1 port map( A => n23317, ZN => n23311);
   U11848 : INV_X1 port map( A => n23317, ZN => n23312);
   U11849 : INV_X1 port map( A => n23316, ZN => n23313);
   U11850 : INV_X1 port map( A => n23294, ZN => n23288);
   U11851 : INV_X1 port map( A => n23294, ZN => n23289);
   U11852 : INV_X1 port map( A => n23293, ZN => n23290);
   U11853 : INV_X1 port map( A => n23656, ZN => n23652);
   U11854 : INV_X1 port map( A => n23596, ZN => n23592);
   U11855 : INV_X1 port map( A => n23616, ZN => n23612);
   U11856 : INV_X1 port map( A => n23636, ZN => n23632);
   U11857 : BUF_X1 port map( A => n23355, Z => n23349);
   U11858 : BUF_X1 port map( A => n23363, Z => n23357);
   U11859 : BUF_X1 port map( A => n23371, Z => n23365);
   U11860 : BUF_X1 port map( A => n23354, Z => n23352);
   U11861 : BUF_X1 port map( A => n23355, Z => n23348);
   U11862 : BUF_X1 port map( A => n23355, Z => n23350);
   U11863 : BUF_X1 port map( A => n23354, Z => n23351);
   U11864 : BUF_X1 port map( A => n23362, Z => n23360);
   U11865 : BUF_X1 port map( A => n23363, Z => n23356);
   U11866 : BUF_X1 port map( A => n23363, Z => n23358);
   U11867 : BUF_X1 port map( A => n23362, Z => n23359);
   U11868 : BUF_X1 port map( A => n23354, Z => n23353);
   U11869 : BUF_X1 port map( A => n23370, Z => n23368);
   U11870 : BUF_X1 port map( A => n23371, Z => n23364);
   U11871 : BUF_X1 port map( A => n23371, Z => n23366);
   U11872 : BUF_X1 port map( A => n23370, Z => n23367);
   U11873 : BUF_X1 port map( A => n23362, Z => n23361);
   U11874 : BUF_X1 port map( A => n23370, Z => n23369);
   U11875 : BUF_X1 port map( A => n23387, Z => n23385);
   U11876 : BUF_X1 port map( A => n23388, Z => n23381);
   U11877 : BUF_X1 port map( A => n23388, Z => n23382);
   U11878 : BUF_X1 port map( A => n23388, Z => n23383);
   U11879 : BUF_X1 port map( A => n23387, Z => n23384);
   U11880 : BUF_X1 port map( A => n23379, Z => n23377);
   U11881 : BUF_X1 port map( A => n23380, Z => n23373);
   U11882 : BUF_X1 port map( A => n23380, Z => n23374);
   U11883 : BUF_X1 port map( A => n23380, Z => n23375);
   U11884 : BUF_X1 port map( A => n23379, Z => n23376);
   U11885 : BUF_X1 port map( A => n23395, Z => n23393);
   U11886 : BUF_X1 port map( A => n23396, Z => n23389);
   U11887 : BUF_X1 port map( A => n23396, Z => n23390);
   U11888 : BUF_X1 port map( A => n23396, Z => n23391);
   U11889 : BUF_X1 port map( A => n23395, Z => n23392);
   U11890 : BUF_X1 port map( A => n23227, Z => n23221);
   U11891 : BUF_X1 port map( A => n23527, Z => n22819);
   U11892 : BUF_X1 port map( A => n23527, Z => n22820);
   U11893 : BUF_X1 port map( A => n23527, Z => n22821);
   U11894 : BUF_X1 port map( A => n23547, Z => n22831);
   U11895 : BUF_X1 port map( A => n23547, Z => n22832);
   U11896 : BUF_X1 port map( A => n23547, Z => n22833);
   U11897 : BUF_X1 port map( A => n23567, Z => n22843);
   U11898 : BUF_X1 port map( A => n23567, Z => n22844);
   U11899 : BUF_X1 port map( A => n23567, Z => n22845);
   U11900 : BUF_X1 port map( A => n23587, Z => n22855);
   U11901 : BUF_X1 port map( A => n23587, Z => n22856);
   U11902 : BUF_X1 port map( A => n23587, Z => n22857);
   U11903 : BUF_X1 port map( A => n23537, Z => n22825);
   U11904 : BUF_X1 port map( A => n23537, Z => n22826);
   U11905 : BUF_X1 port map( A => n23537, Z => n22827);
   U11906 : BUF_X1 port map( A => n23577, Z => n22849);
   U11907 : BUF_X1 port map( A => n23577, Z => n22850);
   U11908 : BUF_X1 port map( A => n23577, Z => n22851);
   U11909 : BUF_X1 port map( A => n23557, Z => n22837);
   U11910 : BUF_X1 port map( A => n23557, Z => n22838);
   U11911 : BUF_X1 port map( A => n23557, Z => n22839);
   U11912 : BUF_X1 port map( A => n23403, Z => n23401);
   U11913 : BUF_X1 port map( A => n23404, Z => n23397);
   U11914 : BUF_X1 port map( A => n23404, Z => n23398);
   U11915 : BUF_X1 port map( A => n23404, Z => n23399);
   U11916 : BUF_X1 port map( A => n23403, Z => n23400);
   U11917 : BUF_X1 port map( A => n23387, Z => n23386);
   U11918 : BUF_X1 port map( A => n23235, Z => n23229);
   U11919 : BUF_X1 port map( A => n23243, Z => n23237);
   U11920 : BUF_X1 port map( A => n23219, Z => n23213);
   U11921 : BUF_X1 port map( A => n23379, Z => n23378);
   U11922 : BUF_X1 port map( A => n23395, Z => n23394);
   U11923 : BUF_X1 port map( A => n23226, Z => n23224);
   U11924 : BUF_X1 port map( A => n23227, Z => n23220);
   U11925 : BUF_X1 port map( A => n23227, Z => n23222);
   U11926 : BUF_X1 port map( A => n23226, Z => n23223);
   U11927 : BUF_X1 port map( A => n23403, Z => n23402);
   U11928 : BUF_X1 port map( A => n23234, Z => n23232);
   U11929 : BUF_X1 port map( A => n23235, Z => n23228);
   U11930 : BUF_X1 port map( A => n23235, Z => n23230);
   U11931 : BUF_X1 port map( A => n23234, Z => n23231);
   U11932 : BUF_X1 port map( A => n23226, Z => n23225);
   U11933 : BUF_X1 port map( A => n23242, Z => n23240);
   U11934 : BUF_X1 port map( A => n23243, Z => n23236);
   U11935 : BUF_X1 port map( A => n23243, Z => n23238);
   U11936 : BUF_X1 port map( A => n23242, Z => n23239);
   U11937 : BUF_X1 port map( A => n23528, Z => n22822);
   U11938 : BUF_X1 port map( A => n23528, Z => n22823);
   U11939 : BUF_X1 port map( A => n23548, Z => n22834);
   U11940 : BUF_X1 port map( A => n23548, Z => n22835);
   U11941 : BUF_X1 port map( A => n23568, Z => n22846);
   U11942 : BUF_X1 port map( A => n23568, Z => n22847);
   U11943 : BUF_X1 port map( A => n23588, Z => n22858);
   U11944 : BUF_X1 port map( A => n23588, Z => n22859);
   U11945 : BUF_X1 port map( A => n23538, Z => n22828);
   U11946 : BUF_X1 port map( A => n23538, Z => n22829);
   U11947 : BUF_X1 port map( A => n23578, Z => n22852);
   U11948 : BUF_X1 port map( A => n23578, Z => n22853);
   U11949 : BUF_X1 port map( A => n23558, Z => n22840);
   U11950 : BUF_X1 port map( A => n23558, Z => n22841);
   U11951 : BUF_X1 port map( A => n23218, Z => n23216);
   U11952 : BUF_X1 port map( A => n23219, Z => n23212);
   U11953 : BUF_X1 port map( A => n23219, Z => n23214);
   U11954 : BUF_X1 port map( A => n23218, Z => n23215);
   U11955 : BUF_X1 port map( A => n23338, Z => n23336);
   U11956 : BUF_X1 port map( A => n23339, Z => n23332);
   U11957 : BUF_X1 port map( A => n23339, Z => n23333);
   U11958 : BUF_X1 port map( A => n23339, Z => n23334);
   U11959 : BUF_X1 port map( A => n23338, Z => n23335);
   U11960 : BUF_X1 port map( A => n23234, Z => n23233);
   U11961 : BUF_X1 port map( A => n23250, Z => n23248);
   U11962 : BUF_X1 port map( A => n23251, Z => n23244);
   U11963 : BUF_X1 port map( A => n23251, Z => n23245);
   U11964 : BUF_X1 port map( A => n23251, Z => n23246);
   U11965 : BUF_X1 port map( A => n23250, Z => n23247);
   U11966 : BUF_X1 port map( A => n23258, Z => n23256);
   U11967 : BUF_X1 port map( A => n23259, Z => n23252);
   U11968 : BUF_X1 port map( A => n23259, Z => n23253);
   U11969 : BUF_X1 port map( A => n23259, Z => n23254);
   U11970 : BUF_X1 port map( A => n23258, Z => n23255);
   U11971 : BUF_X1 port map( A => n23266, Z => n23264);
   U11972 : BUF_X1 port map( A => n23267, Z => n23260);
   U11973 : BUF_X1 port map( A => n23267, Z => n23261);
   U11974 : BUF_X1 port map( A => n23267, Z => n23262);
   U11975 : BUF_X1 port map( A => n23266, Z => n23263);
   U11976 : BUF_X1 port map( A => n23242, Z => n23241);
   U11977 : BUF_X1 port map( A => n23218, Z => n23217);
   U11978 : BUF_X1 port map( A => n23346, Z => n23344);
   U11979 : BUF_X1 port map( A => n23347, Z => n23340);
   U11980 : BUF_X1 port map( A => n23347, Z => n23341);
   U11981 : BUF_X1 port map( A => n23347, Z => n23342);
   U11982 : BUF_X1 port map( A => n23346, Z => n23343);
   U11983 : BUF_X1 port map( A => n23250, Z => n23249);
   U11984 : BUF_X1 port map( A => n23258, Z => n23257);
   U11985 : BUF_X1 port map( A => n23266, Z => n23265);
   U11986 : BUF_X1 port map( A => n23338, Z => n23337);
   U11987 : BUF_X1 port map( A => n23607, Z => n22867);
   U11988 : BUF_X1 port map( A => n23607, Z => n22868);
   U11989 : BUF_X1 port map( A => n23607, Z => n22869);
   U11990 : BUF_X1 port map( A => n23627, Z => n22879);
   U11991 : BUF_X1 port map( A => n23627, Z => n22880);
   U11992 : BUF_X1 port map( A => n23627, Z => n22881);
   U11993 : BUF_X1 port map( A => n23647, Z => n22891);
   U11994 : BUF_X1 port map( A => n23647, Z => n22892);
   U11995 : BUF_X1 port map( A => n23647, Z => n22893);
   U11996 : BUF_X1 port map( A => n23667, Z => n22903);
   U11997 : BUF_X1 port map( A => n23667, Z => n22904);
   U11998 : BUF_X1 port map( A => n23667, Z => n22905);
   U11999 : BUF_X1 port map( A => n23346, Z => n23345);
   U12000 : BUF_X1 port map( A => n23657, Z => n22897);
   U12001 : BUF_X1 port map( A => n23657, Z => n22898);
   U12002 : BUF_X1 port map( A => n23657, Z => n22899);
   U12003 : BUF_X1 port map( A => n23528, Z => n22824);
   U12004 : BUF_X1 port map( A => n23548, Z => n22836);
   U12005 : BUF_X1 port map( A => n23568, Z => n22848);
   U12006 : BUF_X1 port map( A => n23588, Z => n22860);
   U12007 : BUF_X1 port map( A => n23538, Z => n22830);
   U12008 : BUF_X1 port map( A => n23578, Z => n22854);
   U12009 : BUF_X1 port map( A => n23558, Z => n22842);
   U12010 : BUF_X1 port map( A => n23597, Z => n22861);
   U12011 : BUF_X1 port map( A => n23597, Z => n22862);
   U12012 : BUF_X1 port map( A => n23597, Z => n22863);
   U12013 : BUF_X1 port map( A => n23617, Z => n22873);
   U12014 : BUF_X1 port map( A => n23617, Z => n22874);
   U12015 : BUF_X1 port map( A => n23617, Z => n22875);
   U12016 : BUF_X1 port map( A => n23637, Z => n22885);
   U12017 : BUF_X1 port map( A => n23637, Z => n22886);
   U12018 : BUF_X1 port map( A => n23637, Z => n22887);
   U12019 : BUF_X1 port map( A => n23608, Z => n22870);
   U12020 : BUF_X1 port map( A => n23608, Z => n22871);
   U12021 : BUF_X1 port map( A => n23628, Z => n22882);
   U12022 : BUF_X1 port map( A => n23628, Z => n22883);
   U12023 : BUF_X1 port map( A => n23648, Z => n22894);
   U12024 : BUF_X1 port map( A => n23648, Z => n22895);
   U12025 : BUF_X1 port map( A => n23668, Z => n22906);
   U12026 : BUF_X1 port map( A => n23668, Z => n22907);
   U12027 : BUF_X1 port map( A => n23658, Z => n22900);
   U12028 : BUF_X1 port map( A => n23658, Z => n22901);
   U12029 : BUF_X1 port map( A => n23598, Z => n22864);
   U12030 : BUF_X1 port map( A => n23598, Z => n22865);
   U12031 : BUF_X1 port map( A => n23618, Z => n22876);
   U12032 : BUF_X1 port map( A => n23618, Z => n22877);
   U12033 : BUF_X1 port map( A => n23638, Z => n22888);
   U12034 : BUF_X1 port map( A => n23638, Z => n22889);
   U12035 : BUF_X1 port map( A => n23608, Z => n22872);
   U12036 : BUF_X1 port map( A => n23628, Z => n22884);
   U12037 : BUF_X1 port map( A => n23648, Z => n22896);
   U12038 : BUF_X1 port map( A => n23668, Z => n22908);
   U12039 : BUF_X1 port map( A => n23658, Z => n22902);
   U12040 : BUF_X1 port map( A => n23598, Z => n22866);
   U12041 : BUF_X1 port map( A => n23618, Z => n22878);
   U12042 : BUF_X1 port map( A => n23638, Z => n22890);
   U12043 : INV_X1 port map( A => n23413, ZN => n23409);
   U12044 : INV_X1 port map( A => n23413, ZN => n23408);
   U12045 : INV_X1 port map( A => n23479, ZN => n23475);
   U12046 : INV_X1 port map( A => n23479, ZN => n23474);
   U12047 : INV_X1 port map( A => n23466, ZN => n23461);
   U12048 : INV_X1 port map( A => n23424, ZN => n23421);
   U12049 : INV_X1 port map( A => n23424, ZN => n23420);
   U12050 : INV_X1 port map( A => n23412, ZN => n23406);
   U12051 : INV_X1 port map( A => n23466, ZN => n23464);
   U12052 : INV_X1 port map( A => n23467, ZN => n23463);
   U12053 : INV_X1 port map( A => n23467, ZN => n23462);
   U12054 : INV_X1 port map( A => n23412, ZN => n23410);
   U12055 : INV_X1 port map( A => n23412, ZN => n23407);
   U12056 : INV_X1 port map( A => n23478, ZN => n23473);
   U12057 : INV_X1 port map( A => n23477, ZN => n23472);
   U12058 : INV_X1 port map( A => n23423, ZN => n23418);
   U12059 : INV_X1 port map( A => n23423, ZN => n23419);
   U12060 : INV_X1 port map( A => n23425, ZN => n23417);
   U12061 : INV_X1 port map( A => n22989, ZN => n22987);
   U12062 : INV_X1 port map( A => n22992, ZN => n22991);
   U12063 : BUF_X1 port map( A => n23510, Z => n23499);
   U12064 : BUF_X1 port map( A => n23509, Z => n23504);
   U12065 : BUF_X1 port map( A => n23510, Z => n23501);
   U12066 : BUF_X1 port map( A => n23509, Z => n23502);
   U12067 : BUF_X1 port map( A => n23455, Z => n23444);
   U12068 : BUF_X1 port map( A => n23454, Z => n23449);
   U12069 : BUF_X1 port map( A => n23455, Z => n23446);
   U12070 : BUF_X1 port map( A => n23454, Z => n23447);
   U12071 : BUF_X1 port map( A => n23510, Z => n23500);
   U12072 : BUF_X1 port map( A => n23509, Z => n23503);
   U12073 : BUF_X1 port map( A => n23455, Z => n23445);
   U12074 : BUF_X1 port map( A => n23454, Z => n23448);
   U12075 : BUF_X1 port map( A => n23493, Z => n23488);
   U12076 : BUF_X1 port map( A => n23494, Z => n23483);
   U12077 : BUF_X1 port map( A => n23494, Z => n23485);
   U12078 : BUF_X1 port map( A => n23493, Z => n23486);
   U12079 : BUF_X1 port map( A => n23439, Z => n23428);
   U12080 : BUF_X1 port map( A => n23438, Z => n23433);
   U12081 : BUF_X1 port map( A => n23439, Z => n23430);
   U12082 : BUF_X1 port map( A => n23438, Z => n23431);
   U12083 : BUF_X1 port map( A => n23494, Z => n23484);
   U12084 : BUF_X1 port map( A => n23493, Z => n23487);
   U12085 : BUF_X1 port map( A => n23439, Z => n23429);
   U12086 : BUF_X1 port map( A => n23438, Z => n23432);
   U12087 : INV_X1 port map( A => n23520, ZN => n23516);
   U12088 : BUF_X1 port map( A => n23756, Z => n23749);
   U12089 : BUF_X1 port map( A => n23756, Z => n23750);
   U12090 : BUF_X1 port map( A => n23756, Z => n23751);
   U12091 : BUF_X1 port map( A => n23755, Z => n23752);
   U12092 : BUF_X1 port map( A => n23755, Z => n23753);
   U12093 : BUF_X1 port map( A => n23755, Z => n23754);
   U12094 : BUF_X1 port map( A => n22676, Z => n23032);
   U12095 : BUF_X1 port map( A => n23798, Z => n23791);
   U12096 : BUF_X1 port map( A => n23798, Z => n23792);
   U12097 : BUF_X1 port map( A => n23798, Z => n23793);
   U12098 : BUF_X1 port map( A => n23797, Z => n23794);
   U12099 : BUF_X1 port map( A => n23797, Z => n23795);
   U12100 : BUF_X1 port map( A => n23797, Z => n23796);
   U12101 : BUF_X1 port map( A => n23789, Z => n23782);
   U12102 : BUF_X1 port map( A => n23789, Z => n23783);
   U12103 : BUF_X1 port map( A => n23789, Z => n23784);
   U12104 : BUF_X1 port map( A => n23788, Z => n23785);
   U12105 : BUF_X1 port map( A => n23788, Z => n23786);
   U12106 : BUF_X1 port map( A => n23788, Z => n23787);
   U12107 : BUF_X1 port map( A => n23730, Z => n23723);
   U12108 : BUF_X1 port map( A => n23730, Z => n23724);
   U12109 : BUF_X1 port map( A => n23730, Z => n23725);
   U12110 : BUF_X1 port map( A => n23729, Z => n23726);
   U12111 : BUF_X1 port map( A => n23729, Z => n23727);
   U12112 : BUF_X1 port map( A => n23729, Z => n23728);
   U12113 : BUF_X1 port map( A => n23704, Z => n23697);
   U12114 : BUF_X1 port map( A => n23704, Z => n23698);
   U12115 : BUF_X1 port map( A => n23704, Z => n23699);
   U12116 : BUF_X1 port map( A => n23703, Z => n23700);
   U12117 : BUF_X1 port map( A => n23703, Z => n23701);
   U12118 : BUF_X1 port map( A => n23712, Z => n23705);
   U12119 : BUF_X1 port map( A => n23712, Z => n23706);
   U12120 : BUF_X1 port map( A => n23712, Z => n23707);
   U12121 : BUF_X1 port map( A => n23711, Z => n23708);
   U12122 : BUF_X1 port map( A => n23711, Z => n23709);
   U12123 : BUF_X1 port map( A => n23703, Z => n23702);
   U12124 : BUF_X1 port map( A => n23711, Z => n23710);
   U12125 : BUF_X1 port map( A => n23721, Z => n23714);
   U12126 : BUF_X1 port map( A => n23721, Z => n23715);
   U12127 : BUF_X1 port map( A => n23721, Z => n23716);
   U12128 : BUF_X1 port map( A => n23720, Z => n23717);
   U12129 : BUF_X1 port map( A => n23720, Z => n23718);
   U12130 : BUF_X1 port map( A => n23806, Z => n23799);
   U12131 : BUF_X1 port map( A => n23806, Z => n23800);
   U12132 : BUF_X1 port map( A => n23806, Z => n23801);
   U12133 : BUF_X1 port map( A => n23805, Z => n23802);
   U12134 : BUF_X1 port map( A => n23805, Z => n23803);
   U12135 : BUF_X1 port map( A => n23747, Z => n23740);
   U12136 : BUF_X1 port map( A => n23747, Z => n23741);
   U12137 : BUF_X1 port map( A => n23747, Z => n23742);
   U12138 : BUF_X1 port map( A => n23746, Z => n23743);
   U12139 : BUF_X1 port map( A => n23746, Z => n23744);
   U12140 : BUF_X1 port map( A => n23720, Z => n23719);
   U12141 : BUF_X1 port map( A => n23780, Z => n23773);
   U12142 : BUF_X1 port map( A => n23780, Z => n23774);
   U12143 : BUF_X1 port map( A => n23780, Z => n23775);
   U12144 : BUF_X1 port map( A => n23779, Z => n23776);
   U12145 : BUF_X1 port map( A => n23779, Z => n23777);
   U12146 : BUF_X1 port map( A => n23805, Z => n23804);
   U12147 : BUF_X1 port map( A => n23746, Z => n23745);
   U12148 : BUF_X1 port map( A => n23779, Z => n23778);
   U12149 : INV_X1 port map( A => n22998, ZN => n22997);
   U12150 : BUF_X1 port map( A => n23764, Z => n23757);
   U12151 : BUF_X1 port map( A => n23764, Z => n23758);
   U12152 : BUF_X1 port map( A => n23764, Z => n23759);
   U12153 : BUF_X1 port map( A => n23763, Z => n23760);
   U12154 : BUF_X1 port map( A => n23763, Z => n23761);
   U12155 : BUF_X1 port map( A => n23772, Z => n23765);
   U12156 : BUF_X1 port map( A => n23772, Z => n23766);
   U12157 : BUF_X1 port map( A => n23772, Z => n23767);
   U12158 : BUF_X1 port map( A => n23771, Z => n23768);
   U12159 : BUF_X1 port map( A => n23771, Z => n23769);
   U12160 : BUF_X1 port map( A => n23763, Z => n23762);
   U12161 : BUF_X1 port map( A => n23771, Z => n23770);
   U12162 : INV_X1 port map( A => n23525, ZN => n23524);
   U12163 : INV_X1 port map( A => n23525, ZN => n23523);
   U12164 : INV_X1 port map( A => n23545, ZN => n23544);
   U12165 : INV_X1 port map( A => n23545, ZN => n23543);
   U12166 : INV_X1 port map( A => n23565, ZN => n23564);
   U12167 : INV_X1 port map( A => n23565, ZN => n23563);
   U12168 : INV_X1 port map( A => n23585, ZN => n23584);
   U12169 : INV_X1 port map( A => n23585, ZN => n23583);
   U12170 : INV_X1 port map( A => n23535, ZN => n23534);
   U12171 : INV_X1 port map( A => n23535, ZN => n23533);
   U12172 : INV_X1 port map( A => n23575, ZN => n23574);
   U12173 : INV_X1 port map( A => n23575, ZN => n23573);
   U12174 : INV_X1 port map( A => n23555, ZN => n23554);
   U12175 : INV_X1 port map( A => n23555, ZN => n23553);
   U12176 : BUF_X1 port map( A => n23695, Z => n23688);
   U12177 : BUF_X1 port map( A => n23695, Z => n23689);
   U12178 : BUF_X1 port map( A => n23695, Z => n23690);
   U12179 : BUF_X1 port map( A => n23694, Z => n23691);
   U12180 : BUF_X1 port map( A => n23694, Z => n23692);
   U12181 : BUF_X1 port map( A => n23694, Z => n23693);
   U12182 : BUF_X1 port map( A => n23687, Z => n23680);
   U12183 : BUF_X1 port map( A => n23687, Z => n23681);
   U12184 : BUF_X1 port map( A => n23687, Z => n23682);
   U12185 : BUF_X1 port map( A => n23686, Z => n23683);
   U12186 : BUF_X1 port map( A => n23686, Z => n23684);
   U12187 : INV_X1 port map( A => n23327, ZN => n23326);
   U12188 : INV_X1 port map( A => n23304, ZN => n23303);
   U12189 : INV_X1 port map( A => n23327, ZN => n23325);
   U12190 : INV_X1 port map( A => n23304, ZN => n23302);
   U12191 : BUF_X1 port map( A => n23686, Z => n23685);
   U12192 : INV_X1 port map( A => n23315, ZN => n23314);
   U12193 : INV_X1 port map( A => n23292, ZN => n23291);
   U12194 : INV_X1 port map( A => n23605, ZN => n23604);
   U12195 : INV_X1 port map( A => n23605, ZN => n23603);
   U12196 : INV_X1 port map( A => n23625, ZN => n23624);
   U12197 : INV_X1 port map( A => n23625, ZN => n23623);
   U12198 : INV_X1 port map( A => n23645, ZN => n23644);
   U12199 : INV_X1 port map( A => n23645, ZN => n23643);
   U12200 : INV_X1 port map( A => n23665, ZN => n23664);
   U12201 : INV_X1 port map( A => n23665, ZN => n23663);
   U12202 : INV_X1 port map( A => n23655, ZN => n23654);
   U12203 : INV_X1 port map( A => n23655, ZN => n23653);
   U12204 : INV_X1 port map( A => n23595, ZN => n23594);
   U12205 : INV_X1 port map( A => n23595, ZN => n23593);
   U12206 : INV_X1 port map( A => n23615, ZN => n23614);
   U12207 : INV_X1 port map( A => n23615, ZN => n23613);
   U12208 : INV_X1 port map( A => n23635, ZN => n23634);
   U12209 : INV_X1 port map( A => n23635, ZN => n23633);
   U12210 : BUF_X1 port map( A => n23738, Z => n23731);
   U12211 : BUF_X1 port map( A => n23738, Z => n23732);
   U12212 : BUF_X1 port map( A => n23738, Z => n23733);
   U12213 : BUF_X1 port map( A => n23737, Z => n23734);
   U12214 : BUF_X1 port map( A => n23737, Z => n23735);
   U12215 : BUF_X1 port map( A => n23679, Z => n23672);
   U12216 : BUF_X1 port map( A => n23679, Z => n23673);
   U12217 : BUF_X1 port map( A => n23679, Z => n23674);
   U12218 : BUF_X1 port map( A => n23678, Z => n23675);
   U12219 : BUF_X1 port map( A => n23678, Z => n23676);
   U12220 : BUF_X1 port map( A => n23737, Z => n23736);
   U12221 : BUF_X1 port map( A => n23678, Z => n23677);
   U12222 : BUF_X1 port map( A => n23456, Z => n23443);
   U12223 : BUF_X1 port map( A => n23457, Z => n23456);
   U12224 : BUF_X1 port map( A => n23511, Z => n23498);
   U12225 : BUF_X1 port map( A => n23512, Z => n23511);
   U12226 : BUF_X1 port map( A => n23440, Z => n23427);
   U12227 : BUF_X1 port map( A => n23441, Z => n23440);
   U12228 : BUF_X1 port map( A => n23495, Z => n23482);
   U12229 : BUF_X1 port map( A => n23496, Z => n23495);
   U12230 : BUF_X1 port map( A => n23508, Z => n23507);
   U12231 : BUF_X1 port map( A => n23437, Z => n23436);
   U12232 : BUF_X1 port map( A => n23492, Z => n23491);
   U12233 : BUF_X1 port map( A => n23453, Z => n23452);
   U12234 : BUF_X1 port map( A => n23183, Z => n23176);
   U12235 : BUF_X1 port map( A => n23183, Z => n23177);
   U12236 : BUF_X1 port map( A => n23183, Z => n23178);
   U12237 : BUF_X1 port map( A => n23182, Z => n23179);
   U12238 : BUF_X1 port map( A => n23182, Z => n23180);
   U12239 : BUF_X1 port map( A => n22989, Z => n22988);
   U12240 : BUF_X1 port map( A => n23151, Z => n23144);
   U12241 : BUF_X1 port map( A => n23151, Z => n23145);
   U12242 : BUF_X1 port map( A => n23151, Z => n23146);
   U12243 : BUF_X1 port map( A => n23150, Z => n23147);
   U12244 : BUF_X1 port map( A => n23150, Z => n23148);
   U12245 : BUF_X1 port map( A => n23182, Z => n23181);
   U12246 : BUF_X1 port map( A => n23150, Z => n23149);
   U12247 : BUF_X1 port map( A => n22676, Z => n23033);
   U12248 : INV_X1 port map( A => n23465, ZN => n23459);
   U12249 : INV_X1 port map( A => n23465, ZN => n23460);
   U12250 : INV_X1 port map( A => n23411, ZN => n23405);
   U12251 : INV_X1 port map( A => n23476, ZN => n23471);
   U12252 : INV_X1 port map( A => n23422, ZN => n23416);
   U12253 : BUF_X1 port map( A => n23086, Z => n23084);
   U12254 : BUF_X1 port map( A => n23086, Z => n23083);
   U12255 : BUF_X1 port map( A => n23087, Z => n23082);
   U12256 : BUF_X1 port map( A => n23087, Z => n23081);
   U12257 : BUF_X1 port map( A => n23087, Z => n23080);
   U12258 : BUF_X1 port map( A => n23119, Z => n23112);
   U12259 : BUF_X1 port map( A => n23119, Z => n23113);
   U12260 : BUF_X1 port map( A => n23119, Z => n23114);
   U12261 : BUF_X1 port map( A => n23118, Z => n23115);
   U12262 : BUF_X1 port map( A => n23118, Z => n23116);
   U12263 : BUF_X1 port map( A => n23078, Z => n23076);
   U12264 : BUF_X1 port map( A => n23078, Z => n23075);
   U12265 : BUF_X1 port map( A => n23079, Z => n23074);
   U12266 : BUF_X1 port map( A => n23079, Z => n23073);
   U12267 : BUF_X1 port map( A => n23079, Z => n23072);
   U12268 : BUF_X1 port map( A => n23111, Z => n23104);
   U12269 : BUF_X1 port map( A => n23111, Z => n23105);
   U12270 : BUF_X1 port map( A => n23111, Z => n23106);
   U12271 : BUF_X1 port map( A => n23110, Z => n23107);
   U12272 : BUF_X1 port map( A => n23110, Z => n23108);
   U12273 : BUF_X1 port map( A => n23095, Z => n23088);
   U12274 : BUF_X1 port map( A => n23095, Z => n23089);
   U12275 : BUF_X1 port map( A => n23095, Z => n23090);
   U12276 : BUF_X1 port map( A => n23094, Z => n23091);
   U12277 : BUF_X1 port map( A => n23094, Z => n23092);
   U12278 : BUF_X1 port map( A => n23127, Z => n23120);
   U12279 : BUF_X1 port map( A => n23127, Z => n23121);
   U12280 : BUF_X1 port map( A => n23127, Z => n23122);
   U12281 : BUF_X1 port map( A => n23126, Z => n23123);
   U12282 : BUF_X1 port map( A => n23126, Z => n23124);
   U12283 : BUF_X1 port map( A => n23103, Z => n23096);
   U12284 : BUF_X1 port map( A => n23103, Z => n23097);
   U12285 : BUF_X1 port map( A => n23103, Z => n23098);
   U12286 : BUF_X1 port map( A => n23102, Z => n23099);
   U12287 : BUF_X1 port map( A => n23102, Z => n23100);
   U12288 : BUF_X1 port map( A => n23135, Z => n23128);
   U12289 : BUF_X1 port map( A => n23135, Z => n23129);
   U12290 : BUF_X1 port map( A => n23135, Z => n23130);
   U12291 : BUF_X1 port map( A => n23134, Z => n23131);
   U12292 : BUF_X1 port map( A => n23134, Z => n23132);
   U12293 : BUF_X1 port map( A => n23167, Z => n23160);
   U12294 : BUF_X1 port map( A => n23167, Z => n23161);
   U12295 : BUF_X1 port map( A => n23167, Z => n23162);
   U12296 : BUF_X1 port map( A => n23166, Z => n23163);
   U12297 : BUF_X1 port map( A => n23166, Z => n23164);
   U12298 : BUF_X1 port map( A => n23086, Z => n23085);
   U12299 : BUF_X1 port map( A => n23118, Z => n23117);
   U12300 : BUF_X1 port map( A => n23078, Z => n23077);
   U12301 : BUF_X1 port map( A => n23110, Z => n23109);
   U12302 : BUF_X1 port map( A => n23094, Z => n23093);
   U12303 : BUF_X1 port map( A => n23126, Z => n23125);
   U12304 : BUF_X1 port map( A => n23102, Z => n23101);
   U12305 : BUF_X1 port map( A => n23134, Z => n23133);
   U12306 : BUF_X1 port map( A => n23166, Z => n23165);
   U12307 : BUF_X1 port map( A => n23143, Z => n23136);
   U12308 : BUF_X1 port map( A => n23143, Z => n23137);
   U12309 : BUF_X1 port map( A => n23143, Z => n23138);
   U12310 : BUF_X1 port map( A => n23142, Z => n23139);
   U12311 : BUF_X1 port map( A => n23142, Z => n23140);
   U12312 : BUF_X1 port map( A => n23070, Z => n23068);
   U12313 : BUF_X1 port map( A => n23070, Z => n23067);
   U12314 : BUF_X1 port map( A => n23071, Z => n23066);
   U12315 : BUF_X1 port map( A => n23071, Z => n23065);
   U12316 : BUF_X1 port map( A => n23071, Z => n23064);
   U12317 : BUF_X1 port map( A => n23845, Z => n23834);
   U12318 : BUF_X1 port map( A => n23845, Z => n23835);
   U12319 : BUF_X1 port map( A => n23845, Z => n23836);
   U12320 : BUF_X1 port map( A => n23844, Z => n23837);
   U12321 : BUF_X1 port map( A => n23844, Z => n23838);
   U12322 : BUF_X1 port map( A => n23844, Z => n23839);
   U12323 : BUF_X1 port map( A => n23142, Z => n23141);
   U12324 : BUF_X1 port map( A => n23070, Z => n23069);
   U12325 : BUF_X1 port map( A => n23828, Z => n23823);
   U12326 : BUF_X1 port map( A => n23828, Z => n23822);
   U12327 : BUF_X1 port map( A => n23828, Z => n23821);
   U12328 : BUF_X1 port map( A => n23829, Z => n23820);
   U12329 : BUF_X1 port map( A => n23829, Z => n23819);
   U12330 : BUF_X1 port map( A => n23829, Z => n23818);
   U12331 : BUF_X1 port map( A => n23877, Z => n23866);
   U12332 : BUF_X1 port map( A => n23877, Z => n23867);
   U12333 : BUF_X1 port map( A => n23877, Z => n23868);
   U12334 : BUF_X1 port map( A => n23876, Z => n23869);
   U12335 : BUF_X1 port map( A => n23876, Z => n23870);
   U12336 : BUF_X1 port map( A => n23876, Z => n23871);
   U12337 : BUF_X1 port map( A => n23830, Z => n23817);
   U12338 : BUF_X1 port map( A => n23830, Z => n23816);
   U12339 : BUF_X1 port map( A => n23861, Z => n23850);
   U12340 : BUF_X1 port map( A => n23861, Z => n23851);
   U12341 : BUF_X1 port map( A => n23861, Z => n23852);
   U12342 : BUF_X1 port map( A => n23860, Z => n23853);
   U12343 : BUF_X1 port map( A => n23860, Z => n23854);
   U12344 : BUF_X1 port map( A => n23860, Z => n23855);
   U12345 : BUF_X1 port map( A => n23508, Z => n23505);
   U12346 : BUF_X1 port map( A => n23508, Z => n23506);
   U12347 : BUF_X1 port map( A => n23453, Z => n23450);
   U12348 : BUF_X1 port map( A => n23453, Z => n23451);
   U12349 : BUF_X1 port map( A => n23492, Z => n23489);
   U12350 : BUF_X1 port map( A => n23492, Z => n23490);
   U12351 : BUF_X1 port map( A => n23437, Z => n23434);
   U12352 : BUF_X1 port map( A => n23437, Z => n23435);
   U12353 : BUF_X1 port map( A => n22677, Z => n22993);
   U12354 : BUF_X1 port map( A => n24338, Z => n23185);
   U12355 : BUF_X1 port map( A => n24338, Z => n23184);
   U12356 : BUF_X1 port map( A => n24338, Z => n23186);
   U12357 : BUF_X1 port map( A => n24094, Z => n23016);
   U12358 : BUF_X1 port map( A => n24094, Z => n23017);
   U12359 : BUF_X1 port map( A => n24094, Z => n23018);
   U12360 : BUF_X1 port map( A => n23281, Z => n23279);
   U12361 : BUF_X1 port map( A => n23281, Z => n23278);
   U12362 : BUF_X1 port map( A => n23282, Z => n23277);
   U12363 : BUF_X1 port map( A => n23282, Z => n23276);
   U12364 : BUF_X1 port map( A => n23281, Z => n23280);
   U12365 : BUF_X1 port map( A => n23026, Z => n23024);
   U12366 : BUF_X1 port map( A => n23827, Z => n23826);
   U12367 : BUF_X1 port map( A => n23846, Z => n23833);
   U12368 : BUF_X1 port map( A => n23847, Z => n23846);
   U12369 : BUF_X1 port map( A => n23843, Z => n23842);
   U12370 : BUF_X1 port map( A => n23859, Z => n23858);
   U12371 : BUF_X1 port map( A => n23862, Z => n23849);
   U12372 : BUF_X1 port map( A => n23863, Z => n23862);
   U12373 : BUF_X1 port map( A => n23875, Z => n23874);
   U12374 : BUF_X1 port map( A => n23878, Z => n23865);
   U12375 : BUF_X1 port map( A => n23879, Z => n23878);
   U12376 : BUF_X1 port map( A => n23591, Z => n23590);
   U12377 : BUF_X1 port map( A => n23551, Z => n23550);
   U12378 : BUF_X1 port map( A => n23531, Z => n23530);
   U12379 : BUF_X1 port map( A => n23571, Z => n23570);
   U12380 : BUF_X1 port map( A => n23541, Z => n23540);
   U12381 : BUF_X1 port map( A => n23561, Z => n23560);
   U12382 : BUF_X1 port map( A => n23581, Z => n23580);
   U12383 : BUF_X1 port map( A => n22682, Z => n23331);
   U12384 : BUF_X1 port map( A => n22680, Z => n23308);
   U12385 : BUF_X1 port map( A => n22683, Z => n23320);
   U12386 : BUF_X1 port map( A => n22679, Z => n23297);
   U12387 : BUF_X1 port map( A => n23651, Z => n23650);
   U12388 : BUF_X1 port map( A => n23671, Z => n23670);
   U12389 : BUF_X1 port map( A => n23611, Z => n23610);
   U12390 : BUF_X1 port map( A => n23631, Z => n23630);
   U12391 : BUF_X1 port map( A => n23661, Z => n23660);
   U12392 : BUF_X1 port map( A => n23641, Z => n23640);
   U12393 : BUF_X1 port map( A => n23601, Z => n23600);
   U12394 : BUF_X1 port map( A => n23621, Z => n23620);
   U12395 : NAND2_X1 port map( A1 => n21445, A2 => n23498, ZN => n16795);
   U12396 : BUF_X1 port map( A => n22667, Z => n23513);
   U12397 : BUF_X1 port map( A => n22669, Z => n23442);
   U12398 : BUF_X1 port map( A => n22670, Z => n23497);
   U12399 : BUF_X1 port map( A => n22668, Z => n23458);
   U12400 : BUF_X1 port map( A => n22681, Z => n22999);
   U12401 : INV_X1 port map( A => n23981, ZN => n22989);
   U12402 : BUF_X1 port map( A => n23980, Z => n22984);
   U12403 : BUF_X1 port map( A => n23980, Z => n22985);
   U12404 : BUF_X1 port map( A => n23980, Z => n22986);
   U12405 : BUF_X1 port map( A => n23159, Z => n23152);
   U12406 : BUF_X1 port map( A => n23159, Z => n23153);
   U12407 : BUF_X1 port map( A => n23159, Z => n23154);
   U12408 : BUF_X1 port map( A => n23158, Z => n23155);
   U12409 : BUF_X1 port map( A => n23158, Z => n23156);
   U12410 : BUF_X1 port map( A => n23158, Z => n23157);
   U12411 : BUF_X1 port map( A => n23933, Z => n23926);
   U12412 : BUF_X1 port map( A => n23933, Z => n23927);
   U12413 : BUF_X1 port map( A => n23933, Z => n23928);
   U12414 : BUF_X1 port map( A => n23932, Z => n23929);
   U12415 : BUF_X1 port map( A => n23932, Z => n23930);
   U12416 : BUF_X1 port map( A => n23932, Z => n23931);
   U12417 : BUF_X1 port map( A => n22685, Z => n23470);
   U12418 : BUF_X1 port map( A => n22687, Z => n23415);
   U12419 : BUF_X1 port map( A => n22686, Z => n23481);
   U12420 : BUF_X1 port map( A => n22684, Z => n23426);
   U12421 : BUF_X1 port map( A => n23175, Z => n23168);
   U12422 : BUF_X1 port map( A => n23175, Z => n23169);
   U12423 : BUF_X1 port map( A => n23175, Z => n23170);
   U12424 : BUF_X1 port map( A => n23174, Z => n23171);
   U12425 : BUF_X1 port map( A => n23174, Z => n23172);
   U12426 : BUF_X1 port map( A => n23174, Z => n23173);
   U12427 : BUF_X1 port map( A => n23843, Z => n23840);
   U12428 : BUF_X1 port map( A => n23843, Z => n23841);
   U12429 : BUF_X1 port map( A => n23831, Z => n23830);
   U12430 : BUF_X1 port map( A => n23827, Z => n23825);
   U12431 : BUF_X1 port map( A => n23827, Z => n23824);
   U12432 : BUF_X1 port map( A => n23875, Z => n23872);
   U12433 : BUF_X1 port map( A => n23875, Z => n23873);
   U12434 : BUF_X1 port map( A => n23859, Z => n23856);
   U12435 : BUF_X1 port map( A => n23859, Z => n23857);
   U12436 : INV_X1 port map( A => n23273, ZN => n23270);
   U12437 : BUF_X1 port map( A => n23889, Z => n23882);
   U12438 : BUF_X1 port map( A => n23889, Z => n23883);
   U12439 : BUF_X1 port map( A => n23889, Z => n23884);
   U12440 : BUF_X1 port map( A => n23888, Z => n23885);
   U12441 : BUF_X1 port map( A => n23888, Z => n23886);
   U12442 : BUF_X1 port map( A => n23815, Z => n23808);
   U12443 : BUF_X1 port map( A => n23815, Z => n23809);
   U12444 : BUF_X1 port map( A => n23815, Z => n23810);
   U12445 : BUF_X1 port map( A => n23814, Z => n23811);
   U12446 : BUF_X1 port map( A => n23814, Z => n23812);
   U12447 : BUF_X1 port map( A => n23888, Z => n23887);
   U12448 : BUF_X1 port map( A => n23814, Z => n23813);
   U12449 : BUF_X1 port map( A => n23202, Z => n23200);
   U12450 : BUF_X1 port map( A => n23203, Z => n23196);
   U12451 : BUF_X1 port map( A => n23203, Z => n23197);
   U12452 : BUF_X1 port map( A => n23203, Z => n23198);
   U12453 : BUF_X1 port map( A => n23202, Z => n23199);
   U12454 : BUF_X1 port map( A => n23202, Z => n23201);
   U12455 : BUF_X1 port map( A => n23210, Z => n23208);
   U12456 : BUF_X1 port map( A => n23211, Z => n23205);
   U12457 : BUF_X1 port map( A => n23211, Z => n23206);
   U12458 : BUF_X1 port map( A => n23210, Z => n23207);
   U12459 : BUF_X1 port map( A => n23211, Z => n23204);
   U12460 : INV_X1 port map( A => n23271, ZN => n23269);
   U12461 : BUF_X1 port map( A => n23210, Z => n23209);
   U12462 : BUF_X1 port map( A => n23194, Z => n23188);
   U12463 : BUF_X1 port map( A => n23194, Z => n23189);
   U12464 : BUF_X1 port map( A => n23193, Z => n23190);
   U12465 : BUF_X1 port map( A => n23193, Z => n23191);
   U12466 : BUF_X1 port map( A => n23194, Z => n23187);
   U12467 : BUF_X1 port map( A => n23193, Z => n23192);
   U12468 : BUF_X1 port map( A => n23274, Z => n23281);
   U12469 : BUF_X1 port map( A => n23274, Z => n23282);
   U12470 : AND2_X1 port map( A1 => N78, A2 => n22508, ZN => n22678);
   U12471 : INV_X1 port map( A => n16735, ZN => n23521);
   U12472 : BUF_X2 port map( A => n25392, Z => n22946);
   U12473 : BUF_X2 port map( A => n25392, Z => n22943);
   U12474 : BUF_X2 port map( A => n25392, Z => n22945);
   U12475 : BUF_X2 port map( A => n25392, Z => n22944);
   U12476 : CLKBUF_X1 port map( A => n23010, Z => n23008);
   U12477 : INV_X1 port map( A => n22771, ZN => n22776);
   U12478 : AND2_X1 port map( A1 => n16552, A2 => n23826, ZN => n15213);
   U12479 : BUF_X1 port map( A => n21438, Z => n23832);
   U12480 : AND2_X1 port map( A1 => n22693, A2 => n24335, ZN => n22679);
   U12481 : NAND2_X1 port map( A1 => n16552, A2 => n23295, ZN => n15207);
   U12482 : NAND2_X1 port map( A1 => n16552, A2 => n23306, ZN => n15208);
   U12483 : AND2_X1 port map( A1 => n22693, A2 => n24333, ZN => n22680);
   U12484 : NAND2_X1 port map( A1 => n16552, A2 => n23833, ZN => n15217);
   U12485 : BUF_X1 port map( A => n21440, Z => n23848);
   U12486 : AND2_X1 port map( A1 => n23842, A2 => n16555, ZN => n15220);
   U12487 : BUF_X1 port map( A => n21443, Z => n23864);
   U12488 : NAND2_X1 port map( A1 => n23858, A2 => n16555, ZN => n15218);
   U12489 : BUF_X1 port map( A => n21444, Z => n23880);
   U12490 : AND2_X1 port map( A1 => n23874, A2 => n16555, ZN => n15214);
   U12491 : BUF_X1 port map( A => n23054, Z => n23053);
   U12492 : AND3_X1 port map( A1 => n24333, A2 => n24334, A3 => n24332, ZN => 
                           n22682);
   U12493 : AND3_X1 port map( A1 => n24335, A2 => n24334, A3 => n24332, ZN => 
                           n22683);
   U12494 : BUF_X1 port map( A => n22671, Z => n22994);
   U12495 : BUF_X1 port map( A => n21429, Z => n23002);
   U12496 : AND3_X1 port map( A1 => n18526, A2 => n25402, A3 => n25401, ZN => 
                           n22684);
   U12497 : BUF_X1 port map( A => n22671, Z => n22995);
   U12498 : AND3_X1 port map( A1 => n25402, A2 => n18525, A3 => n25400, ZN => 
                           n22685);
   U12499 : AND2_X1 port map( A1 => n23295, A2 => n16555, ZN => n15215);
   U12500 : AND3_X1 port map( A1 => n25402, A2 => n18525, A3 => n18526, ZN => 
                           n22686);
   U12501 : BUF_X1 port map( A => n22671, Z => n22996);
   U12502 : AND2_X1 port map( A1 => n23306, A2 => n16555, ZN => n15223);
   U12503 : AND3_X1 port map( A1 => n25401, A2 => n25402, A3 => n25400, ZN => 
                           n22687);
   U12504 : AND2_X1 port map( A1 => n22498, A2 => n22506, ZN => n22688);
   U12505 : AND2_X1 port map( A1 => n23033, A2 => n24125, ZN => n22689);
   U12506 : CLKBUF_X1 port map( A => n23010, Z => n23007);
   U12507 : INV_X1 port map( A => n16529, ZN => n25407);
   U12508 : BUF_X1 port map( A => n23916, Z => n23909);
   U12509 : INV_X1 port map( A => n22766, ZN => n23945);
   U12510 : BUF_X1 port map( A => n23916, Z => n23910);
   U12511 : BUF_X1 port map( A => n23916, Z => n23911);
   U12512 : BUF_X1 port map( A => n23915, Z => n23912);
   U12513 : BUF_X1 port map( A => n23915, Z => n23913);
   U12514 : BUF_X1 port map( A => n23925, Z => n23918);
   U12515 : BUF_X1 port map( A => n23925, Z => n23919);
   U12516 : BUF_X1 port map( A => n23925, Z => n23920);
   U12517 : BUF_X1 port map( A => n23924, Z => n23921);
   U12518 : BUF_X1 port map( A => n23924, Z => n23922);
   U12519 : BUF_X1 port map( A => n23915, Z => n23914);
   U12520 : BUF_X1 port map( A => n23924, Z => n23923);
   U12521 : BUF_X1 port map( A => n21429, Z => n23001);
   U12522 : BUF_X1 port map( A => n23906, Z => n23899);
   U12523 : BUF_X1 port map( A => n23906, Z => n23900);
   U12524 : BUF_X1 port map( A => n23906, Z => n23901);
   U12525 : BUF_X1 port map( A => n23905, Z => n23902);
   U12526 : BUF_X1 port map( A => n23905, Z => n23903);
   U12527 : BUF_X1 port map( A => n23062, Z => n23060);
   U12528 : BUF_X1 port map( A => n23062, Z => n23059);
   U12529 : BUF_X1 port map( A => n23063, Z => n23058);
   U12530 : BUF_X1 port map( A => n23063, Z => n23057);
   U12531 : BUF_X1 port map( A => n23063, Z => n23056);
   U12532 : BUF_X1 port map( A => n23905, Z => n23904);
   U12533 : BUF_X1 port map( A => n23062, Z => n23061);
   U12534 : BUF_X1 port map( A => n23942, Z => n23935);
   U12535 : BUF_X1 port map( A => n23942, Z => n23936);
   U12536 : BUF_X1 port map( A => n23942, Z => n23937);
   U12537 : BUF_X1 port map( A => n23941, Z => n23938);
   U12538 : BUF_X1 port map( A => n23941, Z => n23939);
   U12539 : BUF_X1 port map( A => n23941, Z => n23940);
   U12540 : BUF_X1 port map( A => n23897, Z => n23890);
   U12541 : BUF_X1 port map( A => n23897, Z => n23891);
   U12542 : BUF_X1 port map( A => n23897, Z => n23892);
   U12543 : BUF_X1 port map( A => n23896, Z => n23893);
   U12544 : BUF_X1 port map( A => n23896, Z => n23894);
   U12545 : BUF_X1 port map( A => n21429, Z => n23000);
   U12546 : BUF_X1 port map( A => n23896, Z => n23895);
   U12547 : AND2_X1 port map( A1 => n23285, A2 => n20834, ZN => n22690);
   U12548 : INV_X1 port map( A => n23946, ZN => n23943);
   U12549 : INV_X1 port map( A => n23946, ZN => n23944);
   U12550 : BUF_X1 port map( A => n23046, Z => n23045);
   U12551 : BUF_X1 port map( A => n23022, Z => n23019);
   U12552 : BUF_X1 port map( A => n23022, Z => n23020);
   U12553 : BUF_X1 port map( A => n23022, Z => n23021);
   U12554 : BUF_X1 port map( A => n23038, Z => n23035);
   U12555 : BUF_X1 port map( A => n23038, Z => n23036);
   U12556 : BUF_X1 port map( A => n23038, Z => n23037);
   U12557 : INV_X1 port map( A => n23005, ZN => n23003);
   U12558 : INV_X1 port map( A => n23005, ZN => n23004);
   U12559 : AOI221_X1 port map( B1 => n22801, B2 => n22036, C1 => n22959, C2 =>
                           n21243, A => n25252, ZN => n25256);
   U12560 : AND2_X1 port map( A1 => n24126, A2 => n24002, ZN => n22691);
   U12561 : BUF_X1 port map( A => n25384, Z => n22948);
   U12562 : BUF_X1 port map( A => n25384, Z => n22950);
   U12563 : BUF_X2 port map( A => n25389, Z => n22953);
   U12564 : BUF_X1 port map( A => n25384, Z => n22949);
   U12565 : BUF_X1 port map( A => n25384, Z => n22930);
   U12566 : BUF_X1 port map( A => n25384, Z => n22931);
   U12567 : BUF_X1 port map( A => n22501, Z => n23274);
   U12568 : BUF_X2 port map( A => n25389, Z => n22952);
   U12569 : BUF_X2 port map( A => n25389, Z => n22954);
   U12570 : BUF_X2 port map( A => n25389, Z => n22955);
   U12571 : BUF_X2 port map( A => n25385, Z => n22976);
   U12572 : BUF_X2 port map( A => n25385, Z => n22978);
   U12573 : BUF_X2 port map( A => n25385, Z => n22979);
   U12574 : BUF_X2 port map( A => n25385, Z => n22977);
   U12575 : XNOR2_X1 port map( A => n24156, B => n24144, ZN => n22692);
   U12576 : NAND4_X1 port map( A1 => n16530, A2 => n16531, A3 => n16532, A4 => 
                           n16533, ZN => n15107);
   U12577 : AOI22_X1 port map( A1 => n23680, A2 => n21972, B1 => n23672, B2 => 
                           n21351, ZN => n16530);
   U12578 : AOI222_X1 port map( A1 => n23705, A2 => n21908, B1 => n23697, B2 =>
                           n21350, C1 => n23688, C2 => n20833, ZN => n16531);
   U12579 : AOI221_X1 port map( B1 => n23740, B2 => n21026, C1 => n23731, C2 =>
                           n21907, A => n16554, ZN => n16532);
   U12580 : NAND4_X1 port map( A1 => n16508, A2 => n16509, A3 => n16510, A4 => 
                           n16511, ZN => n15108);
   U12581 : AOI22_X1 port map( A1 => n23680, A2 => n21973, B1 => n23672, B2 => 
                           n21352, ZN => n16508);
   U12582 : AOI222_X1 port map( A1 => n23705, A2 => n21909, B1 => n23697, B2 =>
                           n21342, C1 => n23688, C2 => n20825, ZN => n16509);
   U12583 : AOI221_X1 port map( B1 => n23740, B2 => n21018, C1 => n23731, C2 =>
                           n21899, A => n16525, ZN => n16510);
   U12584 : NAND4_X1 port map( A1 => n16487, A2 => n16488, A3 => n16489, A4 => 
                           n16490, ZN => n15109);
   U12585 : AOI22_X1 port map( A1 => n23680, A2 => n21974, B1 => n23672, B2 => 
                           n21353, ZN => n16487);
   U12586 : AOI222_X1 port map( A1 => n23705, A2 => n21910, B1 => n23697, B2 =>
                           n21319, C1 => n23688, C2 => n20802, ZN => n16488);
   U12587 : AOI221_X1 port map( B1 => n23740, B2 => n20995, C1 => n23731, C2 =>
                           n21876, A => n16504, ZN => n16489);
   U12588 : NAND4_X1 port map( A1 => n16466, A2 => n16467, A3 => n16468, A4 => 
                           n16469, ZN => n15110);
   U12589 : AOI22_X1 port map( A1 => n23680, A2 => n21975, B1 => n23672, B2 => 
                           n21354, ZN => n16466);
   U12590 : AOI222_X1 port map( A1 => n23705, A2 => n21911, B1 => n23697, B2 =>
                           n21341, C1 => n23688, C2 => n20824, ZN => n16467);
   U12591 : AOI221_X1 port map( B1 => n23740, B2 => n21017, C1 => n23731, C2 =>
                           n21898, A => n16483, ZN => n16468);
   U12592 : NAND4_X1 port map( A1 => n16445, A2 => n16446, A3 => n16447, A4 => 
                           n16448, ZN => n15111);
   U12593 : AOI22_X1 port map( A1 => n23680, A2 => n21976, B1 => n23672, B2 => 
                           n21355, ZN => n16445);
   U12594 : AOI222_X1 port map( A1 => n23705, A2 => n21912, B1 => n23697, B2 =>
                           n21340, C1 => n23688, C2 => n20823, ZN => n16446);
   U12595 : AOI221_X1 port map( B1 => n23740, B2 => n21016, C1 => n23731, C2 =>
                           n21897, A => n16462, ZN => n16447);
   U12596 : NAND4_X1 port map( A1 => n16424, A2 => n16425, A3 => n16426, A4 => 
                           n16427, ZN => n15112);
   U12597 : AOI22_X1 port map( A1 => n23680, A2 => n21977, B1 => n23672, B2 => 
                           n21356, ZN => n16424);
   U12598 : AOI222_X1 port map( A1 => n23705, A2 => n21913, B1 => n23697, B2 =>
                           n21301, C1 => n23688, C2 => n20784, ZN => n16425);
   U12599 : AOI221_X1 port map( B1 => n23740, B2 => n20977, C1 => n23731, C2 =>
                           n21858, A => n16441, ZN => n16426);
   U12600 : NAND4_X1 port map( A1 => n16403, A2 => n16404, A3 => n16405, A4 => 
                           n16406, ZN => n15113);
   U12601 : AOI22_X1 port map( A1 => n23680, A2 => n21978, B1 => n23672, B2 => 
                           n21357, ZN => n16403);
   U12602 : AOI222_X1 port map( A1 => n23705, A2 => n21914, B1 => n23697, B2 =>
                           n21339, C1 => n23688, C2 => n20822, ZN => n16404);
   U12603 : AOI221_X1 port map( B1 => n23740, B2 => n21015, C1 => n23731, C2 =>
                           n21896, A => n16420, ZN => n16405);
   U12604 : NAND4_X1 port map( A1 => n16382, A2 => n16383, A3 => n16384, A4 => 
                           n16385, ZN => n15114);
   U12605 : AOI22_X1 port map( A1 => n23680, A2 => n21979, B1 => n23672, B2 => 
                           n21358, ZN => n16382);
   U12606 : AOI222_X1 port map( A1 => n23705, A2 => n21915, B1 => n23697, B2 =>
                           n21338, C1 => n23688, C2 => n20821, ZN => n16383);
   U12607 : AOI221_X1 port map( B1 => n23740, B2 => n21014, C1 => n23731, C2 =>
                           n21895, A => n16399, ZN => n16384);
   U12608 : NAND4_X1 port map( A1 => n16361, A2 => n16362, A3 => n16363, A4 => 
                           n16364, ZN => n15115);
   U12609 : AOI22_X1 port map( A1 => n23680, A2 => n21980, B1 => n23672, B2 => 
                           n21359, ZN => n16361);
   U12610 : AOI222_X1 port map( A1 => n23705, A2 => n21916, B1 => n23697, B2 =>
                           n21300, C1 => n23688, C2 => n20783, ZN => n16362);
   U12611 : AOI221_X1 port map( B1 => n23740, B2 => n20976, C1 => n23731, C2 =>
                           n21857, A => n16378, ZN => n16363);
   U12612 : NAND4_X1 port map( A1 => n16340, A2 => n16341, A3 => n16342, A4 => 
                           n16343, ZN => n15116);
   U12613 : AOI22_X1 port map( A1 => n23680, A2 => n21981, B1 => n23672, B2 => 
                           n21360, ZN => n16340);
   U12614 : AOI222_X1 port map( A1 => n23705, A2 => n21917, B1 => n23697, B2 =>
                           n21337, C1 => n23688, C2 => n20820, ZN => n16341);
   U12615 : AOI221_X1 port map( B1 => n23740, B2 => n21013, C1 => n23731, C2 =>
                           n21894, A => n16357, ZN => n16342);
   U12616 : NAND4_X1 port map( A1 => n16319, A2 => n16320, A3 => n16321, A4 => 
                           n16322, ZN => n15117);
   U12617 : AOI22_X1 port map( A1 => n23680, A2 => n21982, B1 => n23672, B2 => 
                           n21361, ZN => n16319);
   U12618 : AOI222_X1 port map( A1 => n23705, A2 => n21918, B1 => n23697, B2 =>
                           n21336, C1 => n23688, C2 => n20819, ZN => n16320);
   U12619 : AOI221_X1 port map( B1 => n23740, B2 => n21012, C1 => n23731, C2 =>
                           n21893, A => n16336, ZN => n16321);
   U12620 : NAND4_X1 port map( A1 => n16298, A2 => n16299, A3 => n16300, A4 => 
                           n16301, ZN => n15118);
   U12621 : AOI22_X1 port map( A1 => n23680, A2 => n21983, B1 => n23672, B2 => 
                           n21362, ZN => n16298);
   U12622 : AOI222_X1 port map( A1 => n23705, A2 => n21919, B1 => n23697, B2 =>
                           n21299, C1 => n23688, C2 => n20782, ZN => n16299);
   U12623 : AOI221_X1 port map( B1 => n23740, B2 => n20975, C1 => n23731, C2 =>
                           n21856, A => n16315, ZN => n16300);
   U12624 : NAND4_X1 port map( A1 => n16277, A2 => n16278, A3 => n16279, A4 => 
                           n16280, ZN => n15119);
   U12625 : AOI22_X1 port map( A1 => n23681, A2 => n21984, B1 => n23673, B2 => 
                           n21363, ZN => n16277);
   U12626 : AOI222_X1 port map( A1 => n23706, A2 => n21920, B1 => n23698, B2 =>
                           n21335, C1 => n23689, C2 => n20818, ZN => n16278);
   U12627 : AOI221_X1 port map( B1 => n23741, B2 => n21011, C1 => n23732, C2 =>
                           n21892, A => n16294, ZN => n16279);
   U12628 : NAND4_X1 port map( A1 => n16256, A2 => n16257, A3 => n16258, A4 => 
                           n16259, ZN => n15120);
   U12629 : AOI22_X1 port map( A1 => n23681, A2 => n21985, B1 => n23673, B2 => 
                           n21364, ZN => n16256);
   U12630 : AOI222_X1 port map( A1 => n23706, A2 => n21921, B1 => n23698, B2 =>
                           n21334, C1 => n23689, C2 => n20817, ZN => n16257);
   U12631 : AOI221_X1 port map( B1 => n23741, B2 => n21010, C1 => n23732, C2 =>
                           n21891, A => n16273, ZN => n16258);
   U12632 : NAND4_X1 port map( A1 => n16235, A2 => n16236, A3 => n16237, A4 => 
                           n16238, ZN => n15121);
   U12633 : AOI22_X1 port map( A1 => n23681, A2 => n21986, B1 => n23673, B2 => 
                           n21365, ZN => n16235);
   U12634 : AOI222_X1 port map( A1 => n23706, A2 => n21922, B1 => n23698, B2 =>
                           n21298, C1 => n23689, C2 => n20781, ZN => n16236);
   U12635 : AOI221_X1 port map( B1 => n23741, B2 => n20974, C1 => n23732, C2 =>
                           n21855, A => n16252, ZN => n16237);
   U12636 : NAND4_X1 port map( A1 => n16214, A2 => n16215, A3 => n16216, A4 => 
                           n16217, ZN => n15122);
   U12637 : AOI22_X1 port map( A1 => n23681, A2 => n21987, B1 => n23673, B2 => 
                           n21366, ZN => n16214);
   U12638 : AOI222_X1 port map( A1 => n23706, A2 => n21923, B1 => n23698, B2 =>
                           n21318, C1 => n23689, C2 => n20801, ZN => n16215);
   U12639 : AOI221_X1 port map( B1 => n23741, B2 => n20994, C1 => n23732, C2 =>
                           n21875, A => n16231, ZN => n16216);
   U12640 : NAND4_X1 port map( A1 => n16193, A2 => n16194, A3 => n16195, A4 => 
                           n16196, ZN => n15123);
   U12641 : AOI22_X1 port map( A1 => n23681, A2 => n21988, B1 => n23673, B2 => 
                           n21367, ZN => n16193);
   U12642 : AOI222_X1 port map( A1 => n23706, A2 => n21924, B1 => n23698, B2 =>
                           n21333, C1 => n23689, C2 => n20816, ZN => n16194);
   U12643 : AOI221_X1 port map( B1 => n23741, B2 => n21009, C1 => n23732, C2 =>
                           n21890, A => n16210, ZN => n16195);
   U12644 : NAND4_X1 port map( A1 => n16172, A2 => n16173, A3 => n16174, A4 => 
                           n16175, ZN => n15124);
   U12645 : AOI22_X1 port map( A1 => n23681, A2 => n21989, B1 => n23673, B2 => 
                           n21368, ZN => n16172);
   U12646 : AOI222_X1 port map( A1 => n23706, A2 => n21925, B1 => n23698, B2 =>
                           n21297, C1 => n23689, C2 => n20780, ZN => n16173);
   U12647 : AOI221_X1 port map( B1 => n23741, B2 => n20973, C1 => n23732, C2 =>
                           n21854, A => n16189, ZN => n16174);
   U12648 : NAND4_X1 port map( A1 => n16151, A2 => n16152, A3 => n16153, A4 => 
                           n16154, ZN => n15125);
   U12649 : AOI22_X1 port map( A1 => n23681, A2 => n21990, B1 => n23673, B2 => 
                           n21369, ZN => n16151);
   U12650 : AOI222_X1 port map( A1 => n23706, A2 => n21926, B1 => n23698, B2 =>
                           n21332, C1 => n23689, C2 => n20815, ZN => n16152);
   U12651 : AOI221_X1 port map( B1 => n23741, B2 => n21008, C1 => n23732, C2 =>
                           n21889, A => n16168, ZN => n16153);
   U12652 : NAND4_X1 port map( A1 => n16130, A2 => n16131, A3 => n16132, A4 => 
                           n16133, ZN => n15126);
   U12653 : AOI22_X1 port map( A1 => n23681, A2 => n21991, B1 => n23673, B2 => 
                           n21370, ZN => n16130);
   U12654 : AOI222_X1 port map( A1 => n23706, A2 => n21927, B1 => n23698, B2 =>
                           n21331, C1 => n23689, C2 => n20814, ZN => n16131);
   U12655 : AOI221_X1 port map( B1 => n23741, B2 => n21007, C1 => n23732, C2 =>
                           n21888, A => n16147, ZN => n16132);
   U12656 : NAND4_X1 port map( A1 => n16109, A2 => n16110, A3 => n16111, A4 => 
                           n16112, ZN => n15127);
   U12657 : AOI22_X1 port map( A1 => n23681, A2 => n21992, B1 => n23673, B2 => 
                           n21371, ZN => n16109);
   U12658 : AOI222_X1 port map( A1 => n23706, A2 => n21928, B1 => n23698, B2 =>
                           n21296, C1 => n23689, C2 => n20779, ZN => n16110);
   U12659 : AOI221_X1 port map( B1 => n23741, B2 => n20972, C1 => n23732, C2 =>
                           n21853, A => n16126, ZN => n16111);
   U12660 : NAND4_X1 port map( A1 => n16088, A2 => n16089, A3 => n16090, A4 => 
                           n16091, ZN => n15128);
   U12661 : AOI22_X1 port map( A1 => n23681, A2 => n21993, B1 => n23673, B2 => 
                           n21372, ZN => n16088);
   U12662 : AOI222_X1 port map( A1 => n23706, A2 => n21929, B1 => n23698, B2 =>
                           n21330, C1 => n23689, C2 => n20813, ZN => n16089);
   U12663 : AOI221_X1 port map( B1 => n23741, B2 => n21006, C1 => n23732, C2 =>
                           n21887, A => n16105, ZN => n16090);
   U12664 : NAND4_X1 port map( A1 => n16067, A2 => n16068, A3 => n16069, A4 => 
                           n16070, ZN => n15129);
   U12665 : AOI22_X1 port map( A1 => n23681, A2 => n21994, B1 => n23673, B2 => 
                           n21373, ZN => n16067);
   U12666 : AOI222_X1 port map( A1 => n23706, A2 => n21930, B1 => n23698, B2 =>
                           n21295, C1 => n23689, C2 => n20778, ZN => n16068);
   U12667 : AOI221_X1 port map( B1 => n23741, B2 => n20971, C1 => n23732, C2 =>
                           n21852, A => n16084, ZN => n16069);
   U12668 : NAND4_X1 port map( A1 => n16046, A2 => n16047, A3 => n16048, A4 => 
                           n16049, ZN => n15130);
   U12669 : AOI22_X1 port map( A1 => n23681, A2 => n21995, B1 => n23673, B2 => 
                           n21374, ZN => n16046);
   U12670 : AOI222_X1 port map( A1 => n23706, A2 => n21931, B1 => n23698, B2 =>
                           n21329, C1 => n23689, C2 => n20812, ZN => n16047);
   U12671 : AOI221_X1 port map( B1 => n23741, B2 => n21005, C1 => n23732, C2 =>
                           n21886, A => n16063, ZN => n16048);
   U12672 : NAND4_X1 port map( A1 => n16025, A2 => n16026, A3 => n16027, A4 => 
                           n16028, ZN => n15131);
   U12673 : AOI22_X1 port map( A1 => n23682, A2 => n21996, B1 => n23674, B2 => 
                           n21375, ZN => n16025);
   U12674 : AOI222_X1 port map( A1 => n23707, A2 => n21932, B1 => n23699, B2 =>
                           n21346, C1 => n23690, C2 => n20829, ZN => n16026);
   U12675 : AOI221_X1 port map( B1 => n23742, B2 => n21022, C1 => n23733, C2 =>
                           n21903, A => n16042, ZN => n16027);
   U12676 : NAND4_X1 port map( A1 => n16004, A2 => n16005, A3 => n16006, A4 => 
                           n16007, ZN => n15132);
   U12677 : AOI22_X1 port map( A1 => n23682, A2 => n21997, B1 => n23674, B2 => 
                           n21376, ZN => n16004);
   U12678 : AOI222_X1 port map( A1 => n23707, A2 => n21933, B1 => n23699, B2 =>
                           n21294, C1 => n23690, C2 => n20777, ZN => n16005);
   U12679 : AOI221_X1 port map( B1 => n23742, B2 => n20970, C1 => n23733, C2 =>
                           n21851, A => n16021, ZN => n16006);
   U12680 : NAND4_X1 port map( A1 => n15983, A2 => n15984, A3 => n15985, A4 => 
                           n15986, ZN => n15133);
   U12681 : AOI22_X1 port map( A1 => n23682, A2 => n21998, B1 => n23674, B2 => 
                           n21377, ZN => n15983);
   U12682 : AOI222_X1 port map( A1 => n23707, A2 => n21934, B1 => n23699, B2 =>
                           n21317, C1 => n23690, C2 => n20800, ZN => n15984);
   U12683 : AOI221_X1 port map( B1 => n23742, B2 => n20993, C1 => n23733, C2 =>
                           n21874, A => n16000, ZN => n15985);
   U12684 : NAND4_X1 port map( A1 => n15962, A2 => n15963, A3 => n15964, A4 => 
                           n15965, ZN => n15134);
   U12685 : AOI22_X1 port map( A1 => n23682, A2 => n21999, B1 => n23674, B2 => 
                           n21378, ZN => n15962);
   U12686 : AOI222_X1 port map( A1 => n23707, A2 => n21935, B1 => n23699, B2 =>
                           n21349, C1 => n23690, C2 => n20832, ZN => n15963);
   U12687 : AOI221_X1 port map( B1 => n23742, B2 => n21025, C1 => n23733, C2 =>
                           n21906, A => n15979, ZN => n15964);
   U12688 : NAND4_X1 port map( A1 => n15941, A2 => n15942, A3 => n15943, A4 => 
                           n15944, ZN => n15135);
   U12689 : AOI22_X1 port map( A1 => n23682, A2 => n22000, B1 => n23674, B2 => 
                           n21379, ZN => n15941);
   U12690 : AOI222_X1 port map( A1 => n23707, A2 => n21936, B1 => n23699, B2 =>
                           n21348, C1 => n23690, C2 => n20831, ZN => n15942);
   U12691 : AOI221_X1 port map( B1 => n23742, B2 => n21024, C1 => n23733, C2 =>
                           n21905, A => n15958, ZN => n15943);
   U12692 : NAND4_X1 port map( A1 => n15920, A2 => n15921, A3 => n15922, A4 => 
                           n15923, ZN => n15136);
   U12693 : AOI22_X1 port map( A1 => n23682, A2 => n22001, B1 => n23674, B2 => 
                           n21380, ZN => n15920);
   U12694 : AOI222_X1 port map( A1 => n23707, A2 => n21937, B1 => n23699, B2 =>
                           n21293, C1 => n23690, C2 => n20776, ZN => n15921);
   U12695 : AOI221_X1 port map( B1 => n23742, B2 => n20969, C1 => n23733, C2 =>
                           n21850, A => n15937, ZN => n15922);
   U12696 : NAND4_X1 port map( A1 => n15899, A2 => n15900, A3 => n15901, A4 => 
                           n15902, ZN => n15137);
   U12697 : AOI22_X1 port map( A1 => n23682, A2 => n22002, B1 => n23674, B2 => 
                           n21381, ZN => n15899);
   U12698 : AOI222_X1 port map( A1 => n23707, A2 => n21938, B1 => n23699, B2 =>
                           n21328, C1 => n23690, C2 => n20811, ZN => n15900);
   U12699 : AOI221_X1 port map( B1 => n23742, B2 => n21004, C1 => n23733, C2 =>
                           n21885, A => n15916, ZN => n15901);
   U12700 : NAND4_X1 port map( A1 => n15878, A2 => n15879, A3 => n15880, A4 => 
                           n15881, ZN => n15138);
   U12701 : AOI22_X1 port map( A1 => n23682, A2 => n22003, B1 => n23674, B2 => 
                           n21382, ZN => n15878);
   U12702 : AOI222_X1 port map( A1 => n23707, A2 => n21939, B1 => n23699, B2 =>
                           n21292, C1 => n23690, C2 => n20775, ZN => n15879);
   U12703 : AOI221_X1 port map( B1 => n23742, B2 => n20968, C1 => n23733, C2 =>
                           n21849, A => n15895, ZN => n15880);
   U12704 : NAND4_X1 port map( A1 => n15857, A2 => n15858, A3 => n15859, A4 => 
                           n15860, ZN => n15139);
   U12705 : AOI22_X1 port map( A1 => n23682, A2 => n22004, B1 => n23674, B2 => 
                           n21383, ZN => n15857);
   U12706 : AOI222_X1 port map( A1 => n23707, A2 => n21940, B1 => n23699, B2 =>
                           n21347, C1 => n23690, C2 => n20830, ZN => n15858);
   U12707 : AOI221_X1 port map( B1 => n23742, B2 => n21023, C1 => n23733, C2 =>
                           n21904, A => n15874, ZN => n15859);
   U12708 : NAND4_X1 port map( A1 => n15836, A2 => n15837, A3 => n15838, A4 => 
                           n15839, ZN => n15140);
   U12709 : AOI22_X1 port map( A1 => n23682, A2 => n22005, B1 => n23674, B2 => 
                           n21384, ZN => n15836);
   U12710 : AOI222_X1 port map( A1 => n23707, A2 => n21941, B1 => n23699, B2 =>
                           n21316, C1 => n23690, C2 => n20799, ZN => n15837);
   U12711 : AOI221_X1 port map( B1 => n23742, B2 => n20992, C1 => n23733, C2 =>
                           n21873, A => n15853, ZN => n15838);
   U12712 : NAND4_X1 port map( A1 => n15815, A2 => n15816, A3 => n15817, A4 => 
                           n15818, ZN => n15141);
   U12713 : AOI22_X1 port map( A1 => n23682, A2 => n22006, B1 => n23674, B2 => 
                           n21385, ZN => n15815);
   U12714 : AOI222_X1 port map( A1 => n23707, A2 => n21942, B1 => n23699, B2 =>
                           n21315, C1 => n23690, C2 => n20798, ZN => n15816);
   U12715 : AOI221_X1 port map( B1 => n23742, B2 => n20991, C1 => n23733, C2 =>
                           n21872, A => n15832, ZN => n15817);
   U12716 : NAND4_X1 port map( A1 => n15794, A2 => n15795, A3 => n15796, A4 => 
                           n15797, ZN => n15142);
   U12717 : AOI22_X1 port map( A1 => n23682, A2 => n22007, B1 => n23674, B2 => 
                           n21386, ZN => n15794);
   U12718 : AOI222_X1 port map( A1 => n23707, A2 => n21943, B1 => n23699, B2 =>
                           n21314, C1 => n23690, C2 => n20797, ZN => n15795);
   U12719 : AOI221_X1 port map( B1 => n23742, B2 => n20990, C1 => n23733, C2 =>
                           n21871, A => n15811, ZN => n15796);
   U12720 : NAND4_X1 port map( A1 => n15773, A2 => n15774, A3 => n15775, A4 => 
                           n15776, ZN => n15143);
   U12721 : AOI22_X1 port map( A1 => n23683, A2 => n22008, B1 => n23675, B2 => 
                           n21387, ZN => n15773);
   U12722 : AOI222_X1 port map( A1 => n23708, A2 => n21944, B1 => n23700, B2 =>
                           n21327, C1 => n23691, C2 => n20810, ZN => n15774);
   U12723 : AOI221_X1 port map( B1 => n23743, B2 => n21003, C1 => n23734, C2 =>
                           n21884, A => n15790, ZN => n15775);
   U12724 : NAND4_X1 port map( A1 => n15752, A2 => n15753, A3 => n15754, A4 => 
                           n15755, ZN => n15144);
   U12725 : AOI22_X1 port map( A1 => n23683, A2 => n22009, B1 => n23675, B2 => 
                           n21388, ZN => n15752);
   U12726 : AOI222_X1 port map( A1 => n23708, A2 => n21945, B1 => n23700, B2 =>
                           n21313, C1 => n23691, C2 => n20796, ZN => n15753);
   U12727 : AOI221_X1 port map( B1 => n23743, B2 => n20989, C1 => n23734, C2 =>
                           n21870, A => n15769, ZN => n15754);
   U12728 : NAND4_X1 port map( A1 => n15731, A2 => n15732, A3 => n15733, A4 => 
                           n15734, ZN => n15145);
   U12729 : AOI22_X1 port map( A1 => n23683, A2 => n22010, B1 => n23675, B2 => 
                           n21389, ZN => n15731);
   U12730 : AOI222_X1 port map( A1 => n23708, A2 => n21946, B1 => n23700, B2 =>
                           n21291, C1 => n23691, C2 => n20774, ZN => n15732);
   U12731 : AOI221_X1 port map( B1 => n23743, B2 => n20967, C1 => n23734, C2 =>
                           n21848, A => n15748, ZN => n15733);
   U12732 : NAND4_X1 port map( A1 => n15710, A2 => n15711, A3 => n15712, A4 => 
                           n15713, ZN => n15146);
   U12733 : AOI22_X1 port map( A1 => n23683, A2 => n22011, B1 => n23675, B2 => 
                           n21390, ZN => n15710);
   U12734 : AOI222_X1 port map( A1 => n23708, A2 => n21947, B1 => n23700, B2 =>
                           n21326, C1 => n23691, C2 => n20809, ZN => n15711);
   U12735 : AOI221_X1 port map( B1 => n23743, B2 => n21002, C1 => n23734, C2 =>
                           n21883, A => n15727, ZN => n15712);
   U12736 : NAND4_X1 port map( A1 => n15689, A2 => n15690, A3 => n15691, A4 => 
                           n15692, ZN => n15147);
   U12737 : AOI22_X1 port map( A1 => n23683, A2 => n22012, B1 => n23675, B2 => 
                           n21391, ZN => n15689);
   U12738 : AOI222_X1 port map( A1 => n23708, A2 => n21948, B1 => n23700, B2 =>
                           n21290, C1 => n23691, C2 => n20773, ZN => n15690);
   U12739 : AOI221_X1 port map( B1 => n23743, B2 => n20966, C1 => n23734, C2 =>
                           n21847, A => n15706, ZN => n15691);
   U12740 : NAND4_X1 port map( A1 => n15668, A2 => n15669, A3 => n15670, A4 => 
                           n15671, ZN => n15148);
   U12741 : AOI22_X1 port map( A1 => n23683, A2 => n22013, B1 => n23675, B2 => 
                           n21392, ZN => n15668);
   U12742 : AOI222_X1 port map( A1 => n23708, A2 => n21949, B1 => n23700, B2 =>
                           n21312, C1 => n23691, C2 => n20795, ZN => n15669);
   U12743 : AOI221_X1 port map( B1 => n23743, B2 => n20988, C1 => n23734, C2 =>
                           n21869, A => n15685, ZN => n15670);
   U12744 : NAND4_X1 port map( A1 => n15647, A2 => n15648, A3 => n15649, A4 => 
                           n15650, ZN => n15149);
   U12745 : AOI22_X1 port map( A1 => n23683, A2 => n22014, B1 => n23675, B2 => 
                           n21393, ZN => n15647);
   U12746 : AOI222_X1 port map( A1 => n23708, A2 => n21950, B1 => n23700, B2 =>
                           n21344, C1 => n23691, C2 => n20827, ZN => n15648);
   U12747 : AOI221_X1 port map( B1 => n23743, B2 => n21020, C1 => n23734, C2 =>
                           n21901, A => n15664, ZN => n15649);
   U12748 : NAND4_X1 port map( A1 => n15626, A2 => n15627, A3 => n15628, A4 => 
                           n15629, ZN => n15150);
   U12749 : AOI22_X1 port map( A1 => n23683, A2 => n22015, B1 => n23675, B2 => 
                           n21394, ZN => n15626);
   U12750 : AOI222_X1 port map( A1 => n23708, A2 => n21951, B1 => n23700, B2 =>
                           n21325, C1 => n23691, C2 => n20808, ZN => n15627);
   U12751 : AOI221_X1 port map( B1 => n23743, B2 => n21001, C1 => n23734, C2 =>
                           n21882, A => n15643, ZN => n15628);
   U12752 : NAND4_X1 port map( A1 => n15605, A2 => n15606, A3 => n15607, A4 => 
                           n15608, ZN => n15151);
   U12753 : AOI22_X1 port map( A1 => n23683, A2 => n22016, B1 => n23675, B2 => 
                           n21395, ZN => n15605);
   U12754 : AOI222_X1 port map( A1 => n23708, A2 => n21952, B1 => n23700, B2 =>
                           n21311, C1 => n23691, C2 => n20794, ZN => n15606);
   U12755 : AOI221_X1 port map( B1 => n23743, B2 => n20987, C1 => n23734, C2 =>
                           n21868, A => n15622, ZN => n15607);
   U12756 : NAND4_X1 port map( A1 => n15584, A2 => n15585, A3 => n15586, A4 => 
                           n15587, ZN => n15152);
   U12757 : AOI22_X1 port map( A1 => n23683, A2 => n22017, B1 => n23675, B2 => 
                           n21396, ZN => n15584);
   U12758 : AOI222_X1 port map( A1 => n23708, A2 => n21953, B1 => n23700, B2 =>
                           n21289, C1 => n23691, C2 => n20772, ZN => n15585);
   U12759 : AOI221_X1 port map( B1 => n23743, B2 => n20965, C1 => n23734, C2 =>
                           n21846, A => n15601, ZN => n15586);
   U12760 : NAND4_X1 port map( A1 => n15563, A2 => n15564, A3 => n15565, A4 => 
                           n15566, ZN => n15153);
   U12761 : AOI22_X1 port map( A1 => n23683, A2 => n22018, B1 => n23675, B2 => 
                           n21397, ZN => n15563);
   U12762 : AOI222_X1 port map( A1 => n23708, A2 => n21954, B1 => n23700, B2 =>
                           n21310, C1 => n23691, C2 => n20793, ZN => n15564);
   U12763 : AOI221_X1 port map( B1 => n23743, B2 => n20986, C1 => n23734, C2 =>
                           n21867, A => n15580, ZN => n15565);
   U12764 : NAND4_X1 port map( A1 => n15542, A2 => n15543, A3 => n15544, A4 => 
                           n15545, ZN => n15154);
   U12765 : AOI22_X1 port map( A1 => n23683, A2 => n22019, B1 => n23675, B2 => 
                           n21398, ZN => n15542);
   U12766 : AOI222_X1 port map( A1 => n23708, A2 => n21955, B1 => n23700, B2 =>
                           n21324, C1 => n23691, C2 => n20807, ZN => n15543);
   U12767 : AOI221_X1 port map( B1 => n23743, B2 => n21000, C1 => n23734, C2 =>
                           n21881, A => n15559, ZN => n15544);
   U12768 : NAND4_X1 port map( A1 => n15521, A2 => n15522, A3 => n15523, A4 => 
                           n15524, ZN => n15155);
   U12769 : AOI22_X1 port map( A1 => n23684, A2 => n22020, B1 => n23676, B2 => 
                           n21399, ZN => n15521);
   U12770 : AOI222_X1 port map( A1 => n23709, A2 => n21956, B1 => n23701, B2 =>
                           n21309, C1 => n23692, C2 => n20792, ZN => n15522);
   U12771 : AOI221_X1 port map( B1 => n23744, B2 => n20985, C1 => n23735, C2 =>
                           n21866, A => n15538, ZN => n15523);
   U12772 : NAND4_X1 port map( A1 => n15500, A2 => n15501, A3 => n15502, A4 => 
                           n15503, ZN => n15156);
   U12773 : AOI22_X1 port map( A1 => n23684, A2 => n22021, B1 => n23676, B2 => 
                           n21400, ZN => n15500);
   U12774 : AOI222_X1 port map( A1 => n23709, A2 => n21957, B1 => n23701, B2 =>
                           n21345, C1 => n23692, C2 => n20828, ZN => n15501);
   U12775 : AOI221_X1 port map( B1 => n23744, B2 => n21021, C1 => n23735, C2 =>
                           n21902, A => n15517, ZN => n15502);
   U12776 : NAND4_X1 port map( A1 => n15479, A2 => n15480, A3 => n15481, A4 => 
                           n15482, ZN => n15157);
   U12777 : AOI22_X1 port map( A1 => n23684, A2 => n22022, B1 => n23676, B2 => 
                           n21401, ZN => n15479);
   U12778 : AOI222_X1 port map( A1 => n23709, A2 => n21958, B1 => n23701, B2 =>
                           n21308, C1 => n23692, C2 => n20791, ZN => n15480);
   U12779 : AOI221_X1 port map( B1 => n23744, B2 => n20984, C1 => n23735, C2 =>
                           n21865, A => n15496, ZN => n15481);
   U12780 : NAND4_X1 port map( A1 => n15458, A2 => n15459, A3 => n15460, A4 => 
                           n15461, ZN => n15158);
   U12781 : AOI22_X1 port map( A1 => n23684, A2 => n22023, B1 => n23676, B2 => 
                           n21402, ZN => n15458);
   U12782 : AOI222_X1 port map( A1 => n23709, A2 => n21959, B1 => n23701, B2 =>
                           n21323, C1 => n23692, C2 => n20806, ZN => n15459);
   U12783 : AOI221_X1 port map( B1 => n23744, B2 => n20999, C1 => n23735, C2 =>
                           n21880, A => n15475, ZN => n15460);
   U12784 : NAND4_X1 port map( A1 => n15437, A2 => n15438, A3 => n15439, A4 => 
                           n15440, ZN => n15159);
   U12785 : AOI22_X1 port map( A1 => n23684, A2 => n22024, B1 => n23676, B2 => 
                           n21403, ZN => n15437);
   U12786 : AOI222_X1 port map( A1 => n23709, A2 => n21960, B1 => n23701, B2 =>
                           n21307, C1 => n23692, C2 => n20790, ZN => n15438);
   U12787 : AOI221_X1 port map( B1 => n23744, B2 => n20983, C1 => n23735, C2 =>
                           n21864, A => n15454, ZN => n15439);
   U12788 : NAND4_X1 port map( A1 => n15416, A2 => n15417, A3 => n15418, A4 => 
                           n15419, ZN => n15160);
   U12789 : AOI22_X1 port map( A1 => n23684, A2 => n22025, B1 => n23676, B2 => 
                           n21404, ZN => n15416);
   U12790 : AOI222_X1 port map( A1 => n23709, A2 => n21961, B1 => n23701, B2 =>
                           n21306, C1 => n23692, C2 => n20789, ZN => n15417);
   U12791 : AOI221_X1 port map( B1 => n23744, B2 => n20982, C1 => n23735, C2 =>
                           n21863, A => n15433, ZN => n15418);
   U12792 : NAND4_X1 port map( A1 => n15395, A2 => n15396, A3 => n15397, A4 => 
                           n15398, ZN => n15161);
   U12793 : AOI22_X1 port map( A1 => n23684, A2 => n22026, B1 => n23676, B2 => 
                           n21405, ZN => n15395);
   U12794 : AOI222_X1 port map( A1 => n23709, A2 => n21962, B1 => n23701, B2 =>
                           n21322, C1 => n23692, C2 => n20805, ZN => n15396);
   U12795 : AOI221_X1 port map( B1 => n23744, B2 => n20998, C1 => n23735, C2 =>
                           n21879, A => n15412, ZN => n15397);
   U12796 : NAND4_X1 port map( A1 => n15374, A2 => n15375, A3 => n15376, A4 => 
                           n15377, ZN => n15162);
   U12797 : AOI22_X1 port map( A1 => n23684, A2 => n22027, B1 => n23676, B2 => 
                           n21406, ZN => n15374);
   U12798 : AOI222_X1 port map( A1 => n23709, A2 => n21963, B1 => n23701, B2 =>
                           n21343, C1 => n23692, C2 => n20826, ZN => n15375);
   U12799 : AOI221_X1 port map( B1 => n23744, B2 => n21019, C1 => n23735, C2 =>
                           n21900, A => n15391, ZN => n15376);
   U12800 : NAND4_X1 port map( A1 => n15353, A2 => n15354, A3 => n15355, A4 => 
                           n15356, ZN => n15163);
   U12801 : AOI22_X1 port map( A1 => n23684, A2 => n22028, B1 => n23676, B2 => 
                           n21407, ZN => n15353);
   U12802 : AOI222_X1 port map( A1 => n23709, A2 => n21964, B1 => n23701, B2 =>
                           n21321, C1 => n23692, C2 => n20804, ZN => n15354);
   U12803 : AOI221_X1 port map( B1 => n23744, B2 => n20997, C1 => n23735, C2 =>
                           n21878, A => n15370, ZN => n15355);
   U12804 : NAND4_X1 port map( A1 => n15332, A2 => n15333, A3 => n15334, A4 => 
                           n15335, ZN => n15164);
   U12805 : AOI22_X1 port map( A1 => n23684, A2 => n22029, B1 => n23676, B2 => 
                           n21408, ZN => n15332);
   U12806 : AOI222_X1 port map( A1 => n23709, A2 => n21965, B1 => n23701, B2 =>
                           n21320, C1 => n23692, C2 => n20803, ZN => n15333);
   U12807 : AOI221_X1 port map( B1 => n23744, B2 => n20996, C1 => n23735, C2 =>
                           n21877, A => n15349, ZN => n15334);
   U12808 : NAND4_X1 port map( A1 => n15311, A2 => n15312, A3 => n15313, A4 => 
                           n15314, ZN => n15165);
   U12809 : AOI22_X1 port map( A1 => n23684, A2 => n22030, B1 => n23676, B2 => 
                           n21409, ZN => n15311);
   U12810 : AOI222_X1 port map( A1 => n23709, A2 => n21966, B1 => n23701, B2 =>
                           n21305, C1 => n23692, C2 => n20788, ZN => n15312);
   U12811 : AOI221_X1 port map( B1 => n23744, B2 => n20981, C1 => n23735, C2 =>
                           n21862, A => n15328, ZN => n15313);
   U12812 : NAND4_X1 port map( A1 => n15290, A2 => n15291, A3 => n15292, A4 => 
                           n15293, ZN => n15166);
   U12813 : AOI22_X1 port map( A1 => n23684, A2 => n22031, B1 => n23676, B2 => 
                           n21410, ZN => n15290);
   U12814 : AOI222_X1 port map( A1 => n23709, A2 => n21967, B1 => n23701, B2 =>
                           n21288, C1 => n23692, C2 => n20771, ZN => n15291);
   U12815 : AOI221_X1 port map( B1 => n23744, B2 => n20964, C1 => n23735, C2 =>
                           n21845, A => n15307, ZN => n15292);
   U12816 : NAND4_X1 port map( A1 => n15269, A2 => n15270, A3 => n15271, A4 => 
                           n15272, ZN => n15167);
   U12817 : AOI22_X1 port map( A1 => n23685, A2 => n22032, B1 => n23677, B2 => 
                           n21411, ZN => n15269);
   U12818 : AOI222_X1 port map( A1 => n23710, A2 => n21968, B1 => n23702, B2 =>
                           n21304, C1 => n23693, C2 => n20787, ZN => n15270);
   U12819 : AOI221_X1 port map( B1 => n23745, B2 => n20980, C1 => n23736, C2 =>
                           n21861, A => n15286, ZN => n15271);
   U12820 : NAND4_X1 port map( A1 => n15248, A2 => n15249, A3 => n15250, A4 => 
                           n15251, ZN => n15168);
   U12821 : AOI22_X1 port map( A1 => n23685, A2 => n22033, B1 => n23677, B2 => 
                           n21412, ZN => n15248);
   U12822 : AOI222_X1 port map( A1 => n23710, A2 => n21969, B1 => n23702, B2 =>
                           n21303, C1 => n23693, C2 => n20786, ZN => n15249);
   U12823 : AOI221_X1 port map( B1 => n23745, B2 => n20979, C1 => n23736, C2 =>
                           n21860, A => n15265, ZN => n15250);
   U12824 : NAND4_X1 port map( A1 => n15227, A2 => n15228, A3 => n15229, A4 => 
                           n15230, ZN => n15169);
   U12825 : AOI22_X1 port map( A1 => n23685, A2 => n22034, B1 => n23677, B2 => 
                           n21413, ZN => n15227);
   U12826 : AOI222_X1 port map( A1 => n23710, A2 => n21970, B1 => n23702, B2 =>
                           n21302, C1 => n23693, C2 => n20785, ZN => n15228);
   U12827 : AOI221_X1 port map( B1 => n23745, B2 => n20978, C1 => n23736, C2 =>
                           n21859, A => n15244, ZN => n15229);
   U12828 : NAND4_X1 port map( A1 => n15184, A2 => n15185, A3 => n15186, A4 => 
                           n15187, ZN => n15170);
   U12829 : AOI22_X1 port map( A1 => n23685, A2 => n22035, B1 => n23677, B2 => 
                           n21414, ZN => n15184);
   U12830 : AOI222_X1 port map( A1 => n23710, A2 => n21971, B1 => n23702, B2 =>
                           n21287, C1 => n23693, C2 => n20770, ZN => n15185);
   U12831 : AOI221_X1 port map( B1 => n23745, B2 => n20963, C1 => n23736, C2 =>
                           n21844, A => n15216, ZN => n15186);
   U12832 : AND2_X1 port map( A1 => n24331, A2 => n24336, ZN => n22693);
   U12833 : AND2_X1 port map( A1 => N75, A2 => n23033, ZN => n22694);
   U12834 : BUF_X1 port map( A => n15178, Z => n23934);
   U12835 : NOR3_X1 port map( A1 => n25408, A2 => n25409, A3 => n16529, ZN => 
                           n15178);
   U12836 : NOR2_X1 port map( A1 => n16545, A2 => n16540, ZN => n16552);
   U12837 : NOR2_X1 port map( A1 => n16540, A2 => n25406, ZN => n16555);
   U12838 : AND2_X1 port map( A1 => n24128, A2 => n23036, ZN => n22695);
   U12839 : INV_X1 port map( A => n25394, ZN => n23273);
   U12840 : BUF_X1 port map( A => n15194, Z => n23881);
   U12841 : NAND2_X1 port map( A1 => n25406, A2 => n16540, ZN => n15194);
   U12842 : BUF_X1 port map( A => n15203, Z => n23807);
   U12843 : NAND2_X1 port map( A1 => n16540, A2 => n16545, ZN => n15203);
   U12844 : BUF_X1 port map( A => n25371, Z => n23195);
   U12845 : NOR3_X1 port map( A1 => n16668, A2 => n25404, A3 => n25405, ZN => 
                           n16683);
   U12846 : NAND2_X1 port map( A1 => n25409, A2 => n25408, ZN => n16580);
   U12847 : BUF_X1 port map( A => n25403, Z => n23284);
   U12848 : BUF_X1 port map( A => n25403, Z => n23283);
   U12849 : BUF_X1 port map( A => n23039, Z => n23034);
   U12850 : BUF_X1 port map( A => n24127, Z => n23039);
   U12851 : BUF_X1 port map( A => n25403, Z => n23285);
   U12852 : BUF_X1 port map( A => n22767, Z => n23006);
   U12853 : AND2_X1 port map( A1 => ADD_RD1(2), A2 => n22696, ZN => n22697);
   U12854 : AND2_X1 port map( A1 => n22696, A2 => ADD_RD1(0), ZN => n22698);
   U12855 : NOR2_X1 port map( A1 => n24369, A2 => ADD_RD1(1), ZN => n22699);
   U12856 : NAND3_X1 port map( A1 => n24356, A2 => ADD_RD1(2), A3 => n22484, ZN
                           => n25387);
   U12857 : AND2_X1 port map( A1 => ENABLE, A2 => n5700, ZN => n22700);
   U12858 : OAI22_X1 port map( A1 => n20702, A2 => n23515, B1 => n16635, B2 => 
                           n22815, ZN => n3396);
   U12859 : OAI22_X1 port map( A1 => n20701, A2 => n23515, B1 => n16634, B2 => 
                           n22815, ZN => n3397);
   U12860 : OAI22_X1 port map( A1 => n20700, A2 => n23515, B1 => n16633, B2 => 
                           n22815, ZN => n3398);
   U12861 : OAI22_X1 port map( A1 => n20699, A2 => n23515, B1 => n16632, B2 => 
                           n22815, ZN => n3399);
   U12862 : OAI22_X1 port map( A1 => n20698, A2 => n23515, B1 => n16631, B2 => 
                           n22815, ZN => n3400);
   U12863 : OAI22_X1 port map( A1 => n20697, A2 => n23515, B1 => n16630, B2 => 
                           n22815, ZN => n3401);
   U12864 : OAI22_X1 port map( A1 => n20696, A2 => n23515, B1 => n16629, B2 => 
                           n22818, ZN => n3402);
   U12865 : OAI22_X1 port map( A1 => n20690, A2 => n23514, B1 => n16623, B2 => 
                           n22816, ZN => n3408);
   U12866 : OAI22_X1 port map( A1 => n20689, A2 => n23514, B1 => n16622, B2 => 
                           n22816, ZN => n3409);
   U12867 : OAI22_X1 port map( A1 => n20688, A2 => n23514, B1 => n16621, B2 => 
                           n22816, ZN => n3410);
   U12868 : OAI22_X1 port map( A1 => n20687, A2 => n23514, B1 => n16620, B2 => 
                           n22816, ZN => n3411);
   U12869 : OAI22_X1 port map( A1 => n20686, A2 => n23514, B1 => n16619, B2 => 
                           n22816, ZN => n3412);
   U12870 : OAI22_X1 port map( A1 => n20685, A2 => n23514, B1 => n16618, B2 => 
                           n22816, ZN => n3413);
   U12871 : OAI22_X1 port map( A1 => n20684, A2 => n23514, B1 => n16617, B2 => 
                           n22816, ZN => n3414);
   U12872 : OAI22_X1 port map( A1 => n20678, A2 => n23515, B1 => n16611, B2 => 
                           n22817, ZN => n3420);
   U12873 : OAI22_X1 port map( A1 => n20677, A2 => n23514, B1 => n16610, B2 => 
                           n22817, ZN => n3421);
   U12874 : OAI22_X1 port map( A1 => n20676, A2 => n23516, B1 => n16609, B2 => 
                           n22817, ZN => n3422);
   U12875 : OAI22_X1 port map( A1 => n20675, A2 => n23515, B1 => n16608, B2 => 
                           n22817, ZN => n3423);
   U12876 : OAI22_X1 port map( A1 => n20674, A2 => n23514, B1 => n16607, B2 => 
                           n22817, ZN => n3424);
   U12877 : OAI22_X1 port map( A1 => n20673, A2 => n23516, B1 => n16606, B2 => 
                           n22817, ZN => n3425);
   U12878 : OAI22_X1 port map( A1 => n20672, A2 => n16735, B1 => n16605, B2 => 
                           n22817, ZN => n3426);
   U12879 : OAI22_X1 port map( A1 => n20703, A2 => n23515, B1 => n16636, B2 => 
                           n22815, ZN => n3395);
   U12880 : OAI22_X1 port map( A1 => n20695, A2 => n23515, B1 => n16628, B2 => 
                           n22816, ZN => n3403);
   U12881 : OAI22_X1 port map( A1 => n20694, A2 => n23515, B1 => n16627, B2 => 
                           n22816, ZN => n3404);
   U12882 : OAI22_X1 port map( A1 => n20693, A2 => n23515, B1 => n16626, B2 => 
                           n22816, ZN => n3405);
   U12883 : OAI22_X1 port map( A1 => n20692, A2 => n23515, B1 => n16625, B2 => 
                           n22816, ZN => n3406);
   U12884 : OAI22_X1 port map( A1 => n20691, A2 => n23514, B1 => n16624, B2 => 
                           n22816, ZN => n3407);
   U12885 : OAI22_X1 port map( A1 => n20683, A2 => n23514, B1 => n16616, B2 => 
                           n22817, ZN => n3415);
   U12886 : OAI22_X1 port map( A1 => n20682, A2 => n23514, B1 => n16615, B2 => 
                           n22817, ZN => n3416);
   U12887 : OAI22_X1 port map( A1 => n20681, A2 => n23514, B1 => n16614, B2 => 
                           n22817, ZN => n3417);
   U12888 : OAI22_X1 port map( A1 => n20680, A2 => n23514, B1 => n16613, B2 => 
                           n22817, ZN => n3418);
   U12889 : OAI22_X1 port map( A1 => n20679, A2 => n16735, B1 => n16612, B2 => 
                           n22817, ZN => n3419);
   U12890 : OAI22_X1 port map( A1 => n20671, A2 => n16735, B1 => n16604, B2 => 
                           n22818, ZN => n3427);
   U12891 : OAI22_X1 port map( A1 => n20670, A2 => n16735, B1 => n16603, B2 => 
                           n22818, ZN => n3428);
   U12892 : OAI22_X1 port map( A1 => n20669, A2 => n16735, B1 => n16602, B2 => 
                           n22818, ZN => n3429);
   U12893 : OAI22_X1 port map( A1 => n20668, A2 => n16735, B1 => n16601, B2 => 
                           n22813, ZN => n3430);
   U12894 : OAI22_X1 port map( A1 => n20725, A2 => n23516, B1 => n16658, B2 => 
                           n22813, ZN => n3373);
   U12895 : OAI22_X1 port map( A1 => n20724, A2 => n23516, B1 => n16657, B2 => 
                           n22813, ZN => n3374);
   U12896 : OAI22_X1 port map( A1 => n20723, A2 => n23516, B1 => n16656, B2 => 
                           n22813, ZN => n3375);
   U12897 : OAI22_X1 port map( A1 => n20722, A2 => n23516, B1 => n16655, B2 => 
                           n22813, ZN => n3376);
   U12898 : OAI22_X1 port map( A1 => n20721, A2 => n23516, B1 => n16654, B2 => 
                           n22814, ZN => n3377);
   U12899 : OAI22_X1 port map( A1 => n20720, A2 => n23516, B1 => n16653, B2 => 
                           n22813, ZN => n3378);
   U12900 : OAI22_X1 port map( A1 => n20719, A2 => n23516, B1 => n16652, B2 => 
                           n22814, ZN => n3379);
   U12901 : OAI22_X1 port map( A1 => n20713, A2 => n23516, B1 => n16646, B2 => 
                           n22814, ZN => n3385);
   U12902 : OAI22_X1 port map( A1 => n20712, A2 => n23515, B1 => n16645, B2 => 
                           n22814, ZN => n3386);
   U12903 : OAI22_X1 port map( A1 => n20711, A2 => n23514, B1 => n16644, B2 => 
                           n22814, ZN => n3387);
   U12904 : OAI22_X1 port map( A1 => n20710, A2 => n16735, B1 => n16643, B2 => 
                           n22814, ZN => n3388);
   U12905 : OAI22_X1 port map( A1 => n20709, A2 => n16735, B1 => n16642, B2 => 
                           n22814, ZN => n3389);
   U12906 : OAI22_X1 port map( A1 => n20708, A2 => n16735, B1 => n16641, B2 => 
                           n22814, ZN => n3390);
   U12907 : OAI22_X1 port map( A1 => n20707, A2 => n23516, B1 => n16640, B2 => 
                           n22815, ZN => n3391);
   U12908 : OAI22_X1 port map( A1 => n20727, A2 => n23516, B1 => n16660, B2 => 
                           n22813, ZN => n3371);
   U12909 : OAI22_X1 port map( A1 => n20726, A2 => n23516, B1 => n16659, B2 => 
                           n22813, ZN => n3372);
   U12910 : OAI22_X1 port map( A1 => n20718, A2 => n23516, B1 => n16651, B2 => 
                           n22814, ZN => n3380);
   U12911 : OAI22_X1 port map( A1 => n20717, A2 => n23516, B1 => n16650, B2 => 
                           n22814, ZN => n3381);
   U12912 : OAI22_X1 port map( A1 => n20716, A2 => n23516, B1 => n16649, B2 => 
                           n22814, ZN => n3382);
   U12913 : OAI22_X1 port map( A1 => n20715, A2 => n23515, B1 => n16648, B2 => 
                           n22815, ZN => n3383);
   U12914 : OAI22_X1 port map( A1 => n20714, A2 => n23514, B1 => n16647, B2 => 
                           n22814, ZN => n3384);
   U12915 : OAI22_X1 port map( A1 => n20706, A2 => n23516, B1 => n16639, B2 => 
                           n22815, ZN => n3392);
   U12916 : OAI22_X1 port map( A1 => n20705, A2 => n23515, B1 => n16638, B2 => 
                           n22815, ZN => n3393);
   U12917 : OAI22_X1 port map( A1 => n20704, A2 => n23514, B1 => n16637, B2 => 
                           n22815, ZN => n3394);
   U12918 : OAI22_X1 port map( A1 => n16664, A2 => n22813, B1 => n20731, B2 => 
                           n23516, ZN => n3367);
   U12919 : OAI22_X1 port map( A1 => n20730, A2 => n23516, B1 => n16663, B2 => 
                           n22813, ZN => n3368);
   U12920 : OAI22_X1 port map( A1 => n20729, A2 => n23515, B1 => n16662, B2 => 
                           n22813, ZN => n3369);
   U12921 : OAI22_X1 port map( A1 => n20728, A2 => n23516, B1 => n16661, B2 => 
                           n22813, ZN => n3370);
   U12922 : NOR4_X1 port map( A1 => n16534, A2 => n16535, A3 => n16536, A4 => 
                           n16537, ZN => n16533);
   U12923 : AOI21_X1 port map( B1 => n16543, B2 => n16544, A => n23808, ZN => 
                           n16536);
   U12924 : AOI21_X1 port map( B1 => n16538, B2 => n16539, A => n23882, ZN => 
                           n16537);
   U12925 : OAI22_X1 port map( A1 => n19740, A2 => n23799, B1 => n19804, B2 => 
                           n23791, ZN => n16535);
   U12926 : NOR4_X1 port map( A1 => n16512, A2 => n16513, A3 => n16514, A4 => 
                           n16515, ZN => n16511);
   U12927 : AOI21_X1 port map( B1 => n16520, B2 => n16521, A => n23808, ZN => 
                           n16514);
   U12928 : AOI21_X1 port map( B1 => n16516, B2 => n16517, A => n23882, ZN => 
                           n16515);
   U12929 : OAI22_X1 port map( A1 => n19708, A2 => n23799, B1 => n19772, B2 => 
                           n23791, ZN => n16513);
   U12930 : NOR4_X1 port map( A1 => n16491, A2 => n16492, A3 => n16493, A4 => 
                           n16494, ZN => n16490);
   U12931 : AOI21_X1 port map( B1 => n16499, B2 => n16500, A => n23808, ZN => 
                           n16493);
   U12932 : AOI21_X1 port map( B1 => n16495, B2 => n16496, A => n23882, ZN => 
                           n16494);
   U12933 : OAI22_X1 port map( A1 => n19771, A2 => n23799, B1 => n19835, B2 => 
                           n23791, ZN => n16492);
   U12934 : NOR4_X1 port map( A1 => n16470, A2 => n16471, A3 => n16472, A4 => 
                           n16473, ZN => n16469);
   U12935 : AOI21_X1 port map( B1 => n16478, B2 => n16479, A => n23808, ZN => 
                           n16472);
   U12936 : AOI21_X1 port map( B1 => n16474, B2 => n16475, A => n23882, ZN => 
                           n16473);
   U12937 : OAI22_X1 port map( A1 => n19709, A2 => n23799, B1 => n19773, B2 => 
                           n23791, ZN => n16471);
   U12938 : NOR4_X1 port map( A1 => n16449, A2 => n16450, A3 => n16451, A4 => 
                           n16452, ZN => n16448);
   U12939 : AOI21_X1 port map( B1 => n16457, B2 => n16458, A => n23808, ZN => 
                           n16451);
   U12940 : AOI21_X1 port map( B1 => n16453, B2 => n16454, A => n23882, ZN => 
                           n16452);
   U12941 : OAI22_X1 port map( A1 => n19770, A2 => n23799, B1 => n19834, B2 => 
                           n23791, ZN => n16450);
   U12942 : NOR4_X1 port map( A1 => n16428, A2 => n16429, A3 => n16430, A4 => 
                           n16431, ZN => n16427);
   U12943 : AOI21_X1 port map( B1 => n16436, B2 => n16437, A => n23808, ZN => 
                           n16430);
   U12944 : AOI21_X1 port map( B1 => n16432, B2 => n16433, A => n23882, ZN => 
                           n16431);
   U12945 : OAI22_X1 port map( A1 => n19710, A2 => n23799, B1 => n19774, B2 => 
                           n23791, ZN => n16429);
   U12946 : NOR4_X1 port map( A1 => n16407, A2 => n16408, A3 => n16409, A4 => 
                           n16410, ZN => n16406);
   U12947 : AOI21_X1 port map( B1 => n16415, B2 => n16416, A => n23808, ZN => 
                           n16409);
   U12948 : AOI21_X1 port map( B1 => n16411, B2 => n16412, A => n23882, ZN => 
                           n16410);
   U12949 : OAI22_X1 port map( A1 => n19769, A2 => n23799, B1 => n19833, B2 => 
                           n23791, ZN => n16408);
   U12950 : NOR4_X1 port map( A1 => n16386, A2 => n16387, A3 => n16388, A4 => 
                           n16389, ZN => n16385);
   U12951 : AOI21_X1 port map( B1 => n16394, B2 => n16395, A => n23808, ZN => 
                           n16388);
   U12952 : AOI21_X1 port map( B1 => n16390, B2 => n16391, A => n23882, ZN => 
                           n16389);
   U12953 : OAI22_X1 port map( A1 => n19711, A2 => n23799, B1 => n19775, B2 => 
                           n23791, ZN => n16387);
   U12954 : NOR4_X1 port map( A1 => n16365, A2 => n16366, A3 => n16367, A4 => 
                           n16368, ZN => n16364);
   U12955 : AOI21_X1 port map( B1 => n16373, B2 => n16374, A => n23808, ZN => 
                           n16367);
   U12956 : AOI21_X1 port map( B1 => n16369, B2 => n16370, A => n23882, ZN => 
                           n16368);
   U12957 : OAI22_X1 port map( A1 => n19768, A2 => n23799, B1 => n19832, B2 => 
                           n23791, ZN => n16366);
   U12958 : NOR4_X1 port map( A1 => n16344, A2 => n16345, A3 => n16346, A4 => 
                           n16347, ZN => n16343);
   U12959 : AOI21_X1 port map( B1 => n16352, B2 => n16353, A => n23808, ZN => 
                           n16346);
   U12960 : AOI21_X1 port map( B1 => n16348, B2 => n16349, A => n23882, ZN => 
                           n16347);
   U12961 : OAI22_X1 port map( A1 => n19712, A2 => n23799, B1 => n19776, B2 => 
                           n23791, ZN => n16345);
   U12962 : NOR4_X1 port map( A1 => n16323, A2 => n16324, A3 => n16325, A4 => 
                           n16326, ZN => n16322);
   U12963 : AOI21_X1 port map( B1 => n16331, B2 => n16332, A => n23808, ZN => 
                           n16325);
   U12964 : AOI21_X1 port map( B1 => n16327, B2 => n16328, A => n23882, ZN => 
                           n16326);
   U12965 : OAI22_X1 port map( A1 => n19767, A2 => n23799, B1 => n19831, B2 => 
                           n23791, ZN => n16324);
   U12966 : NOR4_X1 port map( A1 => n16302, A2 => n16303, A3 => n16304, A4 => 
                           n16305, ZN => n16301);
   U12967 : AOI21_X1 port map( B1 => n16310, B2 => n16311, A => n23808, ZN => 
                           n16304);
   U12968 : AOI21_X1 port map( B1 => n16306, B2 => n16307, A => n23882, ZN => 
                           n16305);
   U12969 : OAI22_X1 port map( A1 => n19713, A2 => n23799, B1 => n19777, B2 => 
                           n23791, ZN => n16303);
   U12970 : NOR4_X1 port map( A1 => n16281, A2 => n16282, A3 => n16283, A4 => 
                           n16284, ZN => n16280);
   U12971 : AOI21_X1 port map( B1 => n16289, B2 => n16290, A => n23809, ZN => 
                           n16283);
   U12972 : AOI21_X1 port map( B1 => n16285, B2 => n16286, A => n23883, ZN => 
                           n16284);
   U12973 : OAI22_X1 port map( A1 => n19766, A2 => n23800, B1 => n19830, B2 => 
                           n23792, ZN => n16282);
   U12974 : NOR4_X1 port map( A1 => n16260, A2 => n16261, A3 => n16262, A4 => 
                           n16263, ZN => n16259);
   U12975 : AOI21_X1 port map( B1 => n16268, B2 => n16269, A => n23809, ZN => 
                           n16262);
   U12976 : AOI21_X1 port map( B1 => n16264, B2 => n16265, A => n23883, ZN => 
                           n16263);
   U12977 : OAI22_X1 port map( A1 => n19714, A2 => n23800, B1 => n19778, B2 => 
                           n23792, ZN => n16261);
   U12978 : NOR4_X1 port map( A1 => n16239, A2 => n16240, A3 => n16241, A4 => 
                           n16242, ZN => n16238);
   U12979 : AOI21_X1 port map( B1 => n16247, B2 => n16248, A => n23809, ZN => 
                           n16241);
   U12980 : AOI21_X1 port map( B1 => n16243, B2 => n16244, A => n23883, ZN => 
                           n16242);
   U12981 : OAI22_X1 port map( A1 => n19765, A2 => n23800, B1 => n19829, B2 => 
                           n23792, ZN => n16240);
   U12982 : NOR4_X1 port map( A1 => n16218, A2 => n16219, A3 => n16220, A4 => 
                           n16221, ZN => n16217);
   U12983 : AOI21_X1 port map( B1 => n16226, B2 => n16227, A => n23809, ZN => 
                           n16220);
   U12984 : AOI21_X1 port map( B1 => n16222, B2 => n16223, A => n23883, ZN => 
                           n16221);
   U12985 : OAI22_X1 port map( A1 => n19715, A2 => n23800, B1 => n19779, B2 => 
                           n23792, ZN => n16219);
   U12986 : NOR4_X1 port map( A1 => n16197, A2 => n16198, A3 => n16199, A4 => 
                           n16200, ZN => n16196);
   U12987 : AOI21_X1 port map( B1 => n16205, B2 => n16206, A => n23809, ZN => 
                           n16199);
   U12988 : AOI21_X1 port map( B1 => n16201, B2 => n16202, A => n23883, ZN => 
                           n16200);
   U12989 : OAI22_X1 port map( A1 => n19764, A2 => n23800, B1 => n19828, B2 => 
                           n23792, ZN => n16198);
   U12990 : NOR4_X1 port map( A1 => n16176, A2 => n16177, A3 => n16178, A4 => 
                           n16179, ZN => n16175);
   U12991 : AOI21_X1 port map( B1 => n16184, B2 => n16185, A => n23809, ZN => 
                           n16178);
   U12992 : AOI21_X1 port map( B1 => n16180, B2 => n16181, A => n23883, ZN => 
                           n16179);
   U12993 : OAI22_X1 port map( A1 => n19716, A2 => n23800, B1 => n19780, B2 => 
                           n23792, ZN => n16177);
   U12994 : NOR4_X1 port map( A1 => n16155, A2 => n16156, A3 => n16157, A4 => 
                           n16158, ZN => n16154);
   U12995 : AOI21_X1 port map( B1 => n16163, B2 => n16164, A => n23809, ZN => 
                           n16157);
   U12996 : AOI21_X1 port map( B1 => n16159, B2 => n16160, A => n23883, ZN => 
                           n16158);
   U12997 : OAI22_X1 port map( A1 => n19763, A2 => n23800, B1 => n19827, B2 => 
                           n23792, ZN => n16156);
   U12998 : NOR4_X1 port map( A1 => n16134, A2 => n16135, A3 => n16136, A4 => 
                           n16137, ZN => n16133);
   U12999 : AOI21_X1 port map( B1 => n16142, B2 => n16143, A => n23809, ZN => 
                           n16136);
   U13000 : AOI21_X1 port map( B1 => n16138, B2 => n16139, A => n23883, ZN => 
                           n16137);
   U13001 : OAI22_X1 port map( A1 => n19717, A2 => n23800, B1 => n19781, B2 => 
                           n23792, ZN => n16135);
   U13002 : NOR4_X1 port map( A1 => n16113, A2 => n16114, A3 => n16115, A4 => 
                           n16116, ZN => n16112);
   U13003 : AOI21_X1 port map( B1 => n16121, B2 => n16122, A => n23809, ZN => 
                           n16115);
   U13004 : AOI21_X1 port map( B1 => n16117, B2 => n16118, A => n23883, ZN => 
                           n16116);
   U13005 : OAI22_X1 port map( A1 => n19762, A2 => n23800, B1 => n19826, B2 => 
                           n23792, ZN => n16114);
   U13006 : NOR4_X1 port map( A1 => n16092, A2 => n16093, A3 => n16094, A4 => 
                           n16095, ZN => n16091);
   U13007 : AOI21_X1 port map( B1 => n16100, B2 => n16101, A => n23809, ZN => 
                           n16094);
   U13008 : AOI21_X1 port map( B1 => n16096, B2 => n16097, A => n23883, ZN => 
                           n16095);
   U13009 : OAI22_X1 port map( A1 => n19718, A2 => n23800, B1 => n19782, B2 => 
                           n23792, ZN => n16093);
   U13010 : NOR4_X1 port map( A1 => n16071, A2 => n16072, A3 => n16073, A4 => 
                           n16074, ZN => n16070);
   U13011 : AOI21_X1 port map( B1 => n16079, B2 => n16080, A => n23809, ZN => 
                           n16073);
   U13012 : AOI21_X1 port map( B1 => n16075, B2 => n16076, A => n23883, ZN => 
                           n16074);
   U13013 : OAI22_X1 port map( A1 => n19761, A2 => n23800, B1 => n19825, B2 => 
                           n23792, ZN => n16072);
   U13014 : NOR4_X1 port map( A1 => n16050, A2 => n16051, A3 => n16052, A4 => 
                           n16053, ZN => n16049);
   U13015 : AOI21_X1 port map( B1 => n16058, B2 => n16059, A => n23809, ZN => 
                           n16052);
   U13016 : AOI21_X1 port map( B1 => n16054, B2 => n16055, A => n23883, ZN => 
                           n16053);
   U13017 : OAI22_X1 port map( A1 => n19719, A2 => n23800, B1 => n19783, B2 => 
                           n23792, ZN => n16051);
   U13018 : NOR4_X1 port map( A1 => n16029, A2 => n16030, A3 => n16031, A4 => 
                           n16032, ZN => n16028);
   U13019 : AOI21_X1 port map( B1 => n16037, B2 => n16038, A => n23810, ZN => 
                           n16031);
   U13020 : AOI21_X1 port map( B1 => n16033, B2 => n16034, A => n23884, ZN => 
                           n16032);
   U13021 : OAI22_X1 port map( A1 => n19760, A2 => n23801, B1 => n19824, B2 => 
                           n23793, ZN => n16030);
   U13022 : NOR4_X1 port map( A1 => n16008, A2 => n16009, A3 => n16010, A4 => 
                           n16011, ZN => n16007);
   U13023 : AOI21_X1 port map( B1 => n16016, B2 => n16017, A => n23810, ZN => 
                           n16010);
   U13024 : AOI21_X1 port map( B1 => n16012, B2 => n16013, A => n23884, ZN => 
                           n16011);
   U13025 : OAI22_X1 port map( A1 => n19720, A2 => n23801, B1 => n19784, B2 => 
                           n23793, ZN => n16009);
   U13026 : NOR4_X1 port map( A1 => n15987, A2 => n15988, A3 => n15989, A4 => 
                           n15990, ZN => n15986);
   U13027 : AOI21_X1 port map( B1 => n15995, B2 => n15996, A => n23810, ZN => 
                           n15989);
   U13028 : AOI21_X1 port map( B1 => n15991, B2 => n15992, A => n23884, ZN => 
                           n15990);
   U13029 : OAI22_X1 port map( A1 => n19759, A2 => n23801, B1 => n19823, B2 => 
                           n23793, ZN => n15988);
   U13030 : NOR4_X1 port map( A1 => n15966, A2 => n15967, A3 => n15968, A4 => 
                           n15969, ZN => n15965);
   U13031 : AOI21_X1 port map( B1 => n15974, B2 => n15975, A => n23810, ZN => 
                           n15968);
   U13032 : AOI21_X1 port map( B1 => n15970, B2 => n15971, A => n23884, ZN => 
                           n15969);
   U13033 : OAI22_X1 port map( A1 => n19721, A2 => n23801, B1 => n19785, B2 => 
                           n23793, ZN => n15967);
   U13034 : NOR4_X1 port map( A1 => n15945, A2 => n15946, A3 => n15947, A4 => 
                           n15948, ZN => n15944);
   U13035 : AOI21_X1 port map( B1 => n15953, B2 => n15954, A => n23810, ZN => 
                           n15947);
   U13036 : AOI21_X1 port map( B1 => n15949, B2 => n15950, A => n23884, ZN => 
                           n15948);
   U13037 : OAI22_X1 port map( A1 => n19758, A2 => n23801, B1 => n19822, B2 => 
                           n23793, ZN => n15946);
   U13038 : NOR4_X1 port map( A1 => n15924, A2 => n15925, A3 => n15926, A4 => 
                           n15927, ZN => n15923);
   U13039 : AOI21_X1 port map( B1 => n15932, B2 => n15933, A => n23810, ZN => 
                           n15926);
   U13040 : AOI21_X1 port map( B1 => n15928, B2 => n15929, A => n23884, ZN => 
                           n15927);
   U13041 : OAI22_X1 port map( A1 => n19722, A2 => n23801, B1 => n19786, B2 => 
                           n23793, ZN => n15925);
   U13042 : NOR4_X1 port map( A1 => n15903, A2 => n15904, A3 => n15905, A4 => 
                           n15906, ZN => n15902);
   U13043 : AOI21_X1 port map( B1 => n15911, B2 => n15912, A => n23810, ZN => 
                           n15905);
   U13044 : AOI21_X1 port map( B1 => n15907, B2 => n15908, A => n23884, ZN => 
                           n15906);
   U13045 : OAI22_X1 port map( A1 => n19757, A2 => n23801, B1 => n19821, B2 => 
                           n23793, ZN => n15904);
   U13046 : NOR4_X1 port map( A1 => n15882, A2 => n15883, A3 => n15884, A4 => 
                           n15885, ZN => n15881);
   U13047 : AOI21_X1 port map( B1 => n15890, B2 => n15891, A => n23810, ZN => 
                           n15884);
   U13048 : AOI21_X1 port map( B1 => n15886, B2 => n15887, A => n23884, ZN => 
                           n15885);
   U13049 : OAI22_X1 port map( A1 => n19723, A2 => n23801, B1 => n19787, B2 => 
                           n23793, ZN => n15883);
   U13050 : NOR4_X1 port map( A1 => n15861, A2 => n15862, A3 => n15863, A4 => 
                           n15864, ZN => n15860);
   U13051 : AOI21_X1 port map( B1 => n15869, B2 => n15870, A => n23810, ZN => 
                           n15863);
   U13052 : AOI21_X1 port map( B1 => n15865, B2 => n15866, A => n23884, ZN => 
                           n15864);
   U13053 : OAI22_X1 port map( A1 => n19756, A2 => n23801, B1 => n19820, B2 => 
                           n23793, ZN => n15862);
   U13054 : NOR4_X1 port map( A1 => n15840, A2 => n15841, A3 => n15842, A4 => 
                           n15843, ZN => n15839);
   U13055 : AOI21_X1 port map( B1 => n15848, B2 => n15849, A => n23810, ZN => 
                           n15842);
   U13056 : AOI21_X1 port map( B1 => n15844, B2 => n15845, A => n23884, ZN => 
                           n15843);
   U13057 : OAI22_X1 port map( A1 => n19724, A2 => n23801, B1 => n19788, B2 => 
                           n23793, ZN => n15841);
   U13058 : NOR4_X1 port map( A1 => n15819, A2 => n15820, A3 => n15821, A4 => 
                           n15822, ZN => n15818);
   U13059 : AOI21_X1 port map( B1 => n15827, B2 => n15828, A => n23810, ZN => 
                           n15821);
   U13060 : AOI21_X1 port map( B1 => n15823, B2 => n15824, A => n23884, ZN => 
                           n15822);
   U13061 : OAI22_X1 port map( A1 => n19755, A2 => n23801, B1 => n19819, B2 => 
                           n23793, ZN => n15820);
   U13062 : NOR4_X1 port map( A1 => n15798, A2 => n15799, A3 => n15800, A4 => 
                           n15801, ZN => n15797);
   U13063 : AOI21_X1 port map( B1 => n15806, B2 => n15807, A => n23810, ZN => 
                           n15800);
   U13064 : AOI21_X1 port map( B1 => n15802, B2 => n15803, A => n23884, ZN => 
                           n15801);
   U13065 : OAI22_X1 port map( A1 => n19725, A2 => n23801, B1 => n19789, B2 => 
                           n23793, ZN => n15799);
   U13066 : NOR4_X1 port map( A1 => n15777, A2 => n15778, A3 => n15779, A4 => 
                           n15780, ZN => n15776);
   U13067 : AOI21_X1 port map( B1 => n15785, B2 => n15786, A => n23811, ZN => 
                           n15779);
   U13068 : AOI21_X1 port map( B1 => n15781, B2 => n15782, A => n23885, ZN => 
                           n15780);
   U13069 : OAI22_X1 port map( A1 => n19754, A2 => n23802, B1 => n19818, B2 => 
                           n23794, ZN => n15778);
   U13070 : NOR4_X1 port map( A1 => n15756, A2 => n15757, A3 => n15758, A4 => 
                           n15759, ZN => n15755);
   U13071 : AOI21_X1 port map( B1 => n15764, B2 => n15765, A => n23811, ZN => 
                           n15758);
   U13072 : AOI21_X1 port map( B1 => n15760, B2 => n15761, A => n23885, ZN => 
                           n15759);
   U13073 : OAI22_X1 port map( A1 => n19726, A2 => n23802, B1 => n19790, B2 => 
                           n23794, ZN => n15757);
   U13074 : NOR4_X1 port map( A1 => n15735, A2 => n15736, A3 => n15737, A4 => 
                           n15738, ZN => n15734);
   U13075 : AOI21_X1 port map( B1 => n15743, B2 => n15744, A => n23811, ZN => 
                           n15737);
   U13076 : AOI21_X1 port map( B1 => n15739, B2 => n15740, A => n23885, ZN => 
                           n15738);
   U13077 : OAI22_X1 port map( A1 => n19753, A2 => n23802, B1 => n19817, B2 => 
                           n23794, ZN => n15736);
   U13078 : NOR4_X1 port map( A1 => n15714, A2 => n15715, A3 => n15716, A4 => 
                           n15717, ZN => n15713);
   U13079 : AOI21_X1 port map( B1 => n15722, B2 => n15723, A => n23811, ZN => 
                           n15716);
   U13080 : AOI21_X1 port map( B1 => n15718, B2 => n15719, A => n23885, ZN => 
                           n15717);
   U13081 : OAI22_X1 port map( A1 => n19727, A2 => n23802, B1 => n19791, B2 => 
                           n23794, ZN => n15715);
   U13082 : NOR4_X1 port map( A1 => n15693, A2 => n15694, A3 => n15695, A4 => 
                           n15696, ZN => n15692);
   U13083 : AOI21_X1 port map( B1 => n15701, B2 => n15702, A => n23811, ZN => 
                           n15695);
   U13084 : AOI21_X1 port map( B1 => n15697, B2 => n15698, A => n23885, ZN => 
                           n15696);
   U13085 : OAI22_X1 port map( A1 => n19752, A2 => n23802, B1 => n19816, B2 => 
                           n23794, ZN => n15694);
   U13086 : NOR4_X1 port map( A1 => n15672, A2 => n15673, A3 => n15674, A4 => 
                           n15675, ZN => n15671);
   U13087 : AOI21_X1 port map( B1 => n15680, B2 => n15681, A => n23811, ZN => 
                           n15674);
   U13088 : AOI21_X1 port map( B1 => n15676, B2 => n15677, A => n23885, ZN => 
                           n15675);
   U13089 : OAI22_X1 port map( A1 => n19728, A2 => n23802, B1 => n19792, B2 => 
                           n23794, ZN => n15673);
   U13090 : NOR4_X1 port map( A1 => n15651, A2 => n15652, A3 => n15653, A4 => 
                           n15654, ZN => n15650);
   U13091 : AOI21_X1 port map( B1 => n15659, B2 => n15660, A => n23811, ZN => 
                           n15653);
   U13092 : AOI21_X1 port map( B1 => n15655, B2 => n15656, A => n23885, ZN => 
                           n15654);
   U13093 : OAI22_X1 port map( A1 => n19751, A2 => n23802, B1 => n19815, B2 => 
                           n23794, ZN => n15652);
   U13094 : NOR4_X1 port map( A1 => n15630, A2 => n15631, A3 => n15632, A4 => 
                           n15633, ZN => n15629);
   U13095 : AOI21_X1 port map( B1 => n15638, B2 => n15639, A => n23811, ZN => 
                           n15632);
   U13096 : AOI21_X1 port map( B1 => n15634, B2 => n15635, A => n23885, ZN => 
                           n15633);
   U13097 : OAI22_X1 port map( A1 => n19729, A2 => n23802, B1 => n19793, B2 => 
                           n23794, ZN => n15631);
   U13098 : NOR4_X1 port map( A1 => n15609, A2 => n15610, A3 => n15611, A4 => 
                           n15612, ZN => n15608);
   U13099 : AOI21_X1 port map( B1 => n15617, B2 => n15618, A => n23811, ZN => 
                           n15611);
   U13100 : AOI21_X1 port map( B1 => n15613, B2 => n15614, A => n23885, ZN => 
                           n15612);
   U13101 : OAI22_X1 port map( A1 => n19750, A2 => n23802, B1 => n19814, B2 => 
                           n23794, ZN => n15610);
   U13102 : NOR4_X1 port map( A1 => n15588, A2 => n15589, A3 => n15590, A4 => 
                           n15591, ZN => n15587);
   U13103 : AOI21_X1 port map( B1 => n15596, B2 => n15597, A => n23811, ZN => 
                           n15590);
   U13104 : AOI21_X1 port map( B1 => n15592, B2 => n15593, A => n23885, ZN => 
                           n15591);
   U13105 : OAI22_X1 port map( A1 => n19730, A2 => n23802, B1 => n19794, B2 => 
                           n23794, ZN => n15589);
   U13106 : NOR4_X1 port map( A1 => n15567, A2 => n15568, A3 => n15569, A4 => 
                           n15570, ZN => n15566);
   U13107 : AOI21_X1 port map( B1 => n15575, B2 => n15576, A => n23811, ZN => 
                           n15569);
   U13108 : AOI21_X1 port map( B1 => n15571, B2 => n15572, A => n23885, ZN => 
                           n15570);
   U13109 : OAI22_X1 port map( A1 => n19749, A2 => n23802, B1 => n19813, B2 => 
                           n23794, ZN => n15568);
   U13110 : NOR4_X1 port map( A1 => n15546, A2 => n15547, A3 => n15548, A4 => 
                           n15549, ZN => n15545);
   U13111 : AOI21_X1 port map( B1 => n15554, B2 => n15555, A => n23811, ZN => 
                           n15548);
   U13112 : AOI21_X1 port map( B1 => n15550, B2 => n15551, A => n23885, ZN => 
                           n15549);
   U13113 : OAI22_X1 port map( A1 => n19731, A2 => n23802, B1 => n19795, B2 => 
                           n23794, ZN => n15547);
   U13114 : NOR4_X1 port map( A1 => n15525, A2 => n15526, A3 => n15527, A4 => 
                           n15528, ZN => n15524);
   U13115 : AOI21_X1 port map( B1 => n15533, B2 => n15534, A => n23812, ZN => 
                           n15527);
   U13116 : AOI21_X1 port map( B1 => n15529, B2 => n15530, A => n23886, ZN => 
                           n15528);
   U13117 : OAI22_X1 port map( A1 => n19748, A2 => n23803, B1 => n19812, B2 => 
                           n23795, ZN => n15526);
   U13118 : NOR4_X1 port map( A1 => n15504, A2 => n15505, A3 => n15506, A4 => 
                           n15507, ZN => n15503);
   U13119 : AOI21_X1 port map( B1 => n15512, B2 => n15513, A => n23812, ZN => 
                           n15506);
   U13120 : AOI21_X1 port map( B1 => n15508, B2 => n15509, A => n23886, ZN => 
                           n15507);
   U13121 : OAI22_X1 port map( A1 => n19732, A2 => n23803, B1 => n19796, B2 => 
                           n23795, ZN => n15505);
   U13122 : NOR4_X1 port map( A1 => n15483, A2 => n15484, A3 => n15485, A4 => 
                           n15486, ZN => n15482);
   U13123 : AOI21_X1 port map( B1 => n15491, B2 => n15492, A => n23812, ZN => 
                           n15485);
   U13124 : AOI21_X1 port map( B1 => n15487, B2 => n15488, A => n23886, ZN => 
                           n15486);
   U13125 : OAI22_X1 port map( A1 => n19747, A2 => n23803, B1 => n19811, B2 => 
                           n23795, ZN => n15484);
   U13126 : NOR4_X1 port map( A1 => n15462, A2 => n15463, A3 => n15464, A4 => 
                           n15465, ZN => n15461);
   U13127 : AOI21_X1 port map( B1 => n15470, B2 => n15471, A => n23812, ZN => 
                           n15464);
   U13128 : AOI21_X1 port map( B1 => n15466, B2 => n15467, A => n23886, ZN => 
                           n15465);
   U13129 : OAI22_X1 port map( A1 => n19733, A2 => n23803, B1 => n19797, B2 => 
                           n23795, ZN => n15463);
   U13130 : NOR4_X1 port map( A1 => n15441, A2 => n15442, A3 => n15443, A4 => 
                           n15444, ZN => n15440);
   U13131 : AOI21_X1 port map( B1 => n15449, B2 => n15450, A => n23812, ZN => 
                           n15443);
   U13132 : AOI21_X1 port map( B1 => n15445, B2 => n15446, A => n23886, ZN => 
                           n15444);
   U13133 : OAI22_X1 port map( A1 => n19746, A2 => n23803, B1 => n19810, B2 => 
                           n23795, ZN => n15442);
   U13134 : NOR4_X1 port map( A1 => n15420, A2 => n15421, A3 => n15422, A4 => 
                           n15423, ZN => n15419);
   U13135 : AOI21_X1 port map( B1 => n15428, B2 => n15429, A => n23812, ZN => 
                           n15422);
   U13136 : AOI21_X1 port map( B1 => n15424, B2 => n15425, A => n23886, ZN => 
                           n15423);
   U13137 : OAI22_X1 port map( A1 => n19734, A2 => n23803, B1 => n19798, B2 => 
                           n23795, ZN => n15421);
   U13138 : NOR4_X1 port map( A1 => n15399, A2 => n15400, A3 => n15401, A4 => 
                           n15402, ZN => n15398);
   U13139 : AOI21_X1 port map( B1 => n15407, B2 => n15408, A => n23812, ZN => 
                           n15401);
   U13140 : AOI21_X1 port map( B1 => n15403, B2 => n15404, A => n23886, ZN => 
                           n15402);
   U13141 : OAI22_X1 port map( A1 => n19745, A2 => n23803, B1 => n19809, B2 => 
                           n23795, ZN => n15400);
   U13142 : NOR4_X1 port map( A1 => n15378, A2 => n15379, A3 => n15380, A4 => 
                           n15381, ZN => n15377);
   U13143 : AOI21_X1 port map( B1 => n15386, B2 => n15387, A => n23812, ZN => 
                           n15380);
   U13144 : AOI21_X1 port map( B1 => n15382, B2 => n15383, A => n23886, ZN => 
                           n15381);
   U13145 : OAI22_X1 port map( A1 => n19735, A2 => n23803, B1 => n19799, B2 => 
                           n23795, ZN => n15379);
   U13146 : NOR4_X1 port map( A1 => n15357, A2 => n15358, A3 => n15359, A4 => 
                           n15360, ZN => n15356);
   U13147 : AOI21_X1 port map( B1 => n15365, B2 => n15366, A => n23812, ZN => 
                           n15359);
   U13148 : AOI21_X1 port map( B1 => n15361, B2 => n15362, A => n23886, ZN => 
                           n15360);
   U13149 : OAI22_X1 port map( A1 => n19744, A2 => n23803, B1 => n19808, B2 => 
                           n23795, ZN => n15358);
   U13150 : NOR4_X1 port map( A1 => n15336, A2 => n15337, A3 => n15338, A4 => 
                           n15339, ZN => n15335);
   U13151 : AOI21_X1 port map( B1 => n15344, B2 => n15345, A => n23812, ZN => 
                           n15338);
   U13152 : AOI21_X1 port map( B1 => n15340, B2 => n15341, A => n23886, ZN => 
                           n15339);
   U13153 : OAI22_X1 port map( A1 => n19736, A2 => n23803, B1 => n19800, B2 => 
                           n23795, ZN => n15337);
   U13154 : NOR4_X1 port map( A1 => n15315, A2 => n15316, A3 => n15317, A4 => 
                           n15318, ZN => n15314);
   U13155 : AOI21_X1 port map( B1 => n15323, B2 => n15324, A => n23812, ZN => 
                           n15317);
   U13156 : AOI21_X1 port map( B1 => n15319, B2 => n15320, A => n23886, ZN => 
                           n15318);
   U13157 : OAI22_X1 port map( A1 => n19743, A2 => n23803, B1 => n19807, B2 => 
                           n23795, ZN => n15316);
   U13158 : NOR4_X1 port map( A1 => n15294, A2 => n15295, A3 => n15296, A4 => 
                           n15297, ZN => n15293);
   U13159 : AOI21_X1 port map( B1 => n15302, B2 => n15303, A => n23812, ZN => 
                           n15296);
   U13160 : AOI21_X1 port map( B1 => n15298, B2 => n15299, A => n23886, ZN => 
                           n15297);
   U13161 : OAI22_X1 port map( A1 => n19737, A2 => n23803, B1 => n19801, B2 => 
                           n23795, ZN => n15295);
   U13162 : OAI221_X1 port map( B1 => n19932, B2 => n23782, C1 => n19868, C2 =>
                           n23773, A => n16553, ZN => n16534);
   U13163 : AOI222_X1 port map( A1 => n23765, A2 => n21763, B1 => n23757, B2 =>
                           n21272, C1 => n23749, C2 => n20898, ZN => n16553);
   U13164 : OAI221_X1 port map( B1 => n19900, B2 => n23782, C1 => n19836, C2 =>
                           n23773, A => n16524, ZN => n16512);
   U13165 : AOI222_X1 port map( A1 => n23765, A2 => n21515, B1 => n23757, B2 =>
                           n21086, C1 => n23749, C2 => n20890, ZN => n16524);
   U13166 : OAI221_X1 port map( B1 => n19963, B2 => n23782, C1 => n19899, C2 =>
                           n23773, A => n16503, ZN => n16491);
   U13167 : AOI222_X1 port map( A1 => n23765, A2 => n21512, B1 => n23757, B2 =>
                           n21083, C1 => n23749, C2 => n20887, ZN => n16503);
   U13168 : OAI221_X1 port map( B1 => n19901, B2 => n23782, C1 => n19837, C2 =>
                           n23773, A => n16482, ZN => n16470);
   U13169 : AOI222_X1 port map( A1 => n23765, A2 => n21514, B1 => n23757, B2 =>
                           n21085, C1 => n23749, C2 => n20889, ZN => n16482);
   U13170 : OAI221_X1 port map( B1 => n19962, B2 => n23782, C1 => n19898, C2 =>
                           n23773, A => n16461, ZN => n16449);
   U13171 : AOI222_X1 port map( A1 => n23765, A2 => n21513, B1 => n23757, B2 =>
                           n21084, C1 => n23749, C2 => n20888, ZN => n16461);
   U13172 : OAI221_X1 port map( B1 => n19902, B2 => n23782, C1 => n19838, C2 =>
                           n23773, A => n16440, ZN => n16428);
   U13173 : AOI222_X1 port map( A1 => n23765, A2 => n21471, B1 => n23757, B2 =>
                           n21042, C1 => n23749, C2 => n20846, ZN => n16440);
   U13174 : OAI221_X1 port map( B1 => n19961, B2 => n23782, C1 => n19897, C2 =>
                           n23773, A => n16419, ZN => n16407);
   U13175 : AOI222_X1 port map( A1 => n23765, A2 => n21501, B1 => n23757, B2 =>
                           n21072, C1 => n23749, C2 => n20876, ZN => n16419);
   U13176 : OAI221_X1 port map( B1 => n19903, B2 => n23782, C1 => n19839, C2 =>
                           n23773, A => n16398, ZN => n16386);
   U13177 : AOI222_X1 port map( A1 => n23765, A2 => n21498, B1 => n23757, B2 =>
                           n21069, C1 => n23749, C2 => n20873, ZN => n16398);
   U13178 : OAI221_X1 port map( B1 => n19960, B2 => n23782, C1 => n19896, C2 =>
                           n23773, A => n16377, ZN => n16365);
   U13179 : AOI222_X1 port map( A1 => n23765, A2 => n21463, B1 => n23757, B2 =>
                           n21034, C1 => n23749, C2 => n20838, ZN => n16377);
   U13180 : OAI221_X1 port map( B1 => n19904, B2 => n23782, C1 => n19840, C2 =>
                           n23773, A => n16356, ZN => n16344);
   U13181 : AOI222_X1 port map( A1 => n23765, A2 => n21497, B1 => n23757, B2 =>
                           n21068, C1 => n23749, C2 => n20872, ZN => n16356);
   U13182 : OAI221_X1 port map( B1 => n19959, B2 => n23782, C1 => n19895, C2 =>
                           n23773, A => n16335, ZN => n16323);
   U13183 : AOI222_X1 port map( A1 => n23765, A2 => n21499, B1 => n23757, B2 =>
                           n21070, C1 => n23749, C2 => n20874, ZN => n16335);
   U13184 : OAI221_X1 port map( B1 => n19905, B2 => n23782, C1 => n19841, C2 =>
                           n23773, A => n16314, ZN => n16302);
   U13185 : AOI222_X1 port map( A1 => n23765, A2 => n21466, B1 => n23757, B2 =>
                           n21037, C1 => n23749, C2 => n20841, ZN => n16314);
   U13186 : OAI221_X1 port map( B1 => n19958, B2 => n23783, C1 => n19894, C2 =>
                           n23774, A => n16293, ZN => n16281);
   U13187 : AOI222_X1 port map( A1 => n23766, A2 => n21505, B1 => n23758, B2 =>
                           n21076, C1 => n23750, C2 => n20880, ZN => n16293);
   U13188 : OAI221_X1 port map( B1 => n19906, B2 => n23783, C1 => n19842, C2 =>
                           n23774, A => n16272, ZN => n16260);
   U13189 : AOI222_X1 port map( A1 => n23766, A2 => n21496, B1 => n23758, B2 =>
                           n21067, C1 => n23750, C2 => n20871, ZN => n16272);
   U13190 : OAI221_X1 port map( B1 => n19957, B2 => n23783, C1 => n19893, C2 =>
                           n23774, A => n16251, ZN => n16239);
   U13191 : AOI222_X1 port map( A1 => n23766, A2 => n21470, B1 => n23758, B2 =>
                           n21041, C1 => n23750, C2 => n20845, ZN => n16251);
   U13192 : OAI221_X1 port map( B1 => n19907, B2 => n23783, C1 => n19843, C2 =>
                           n23774, A => n16230, ZN => n16218);
   U13193 : AOI222_X1 port map( A1 => n23766, A2 => n21489, B1 => n23758, B2 =>
                           n21060, C1 => n23750, C2 => n20864, ZN => n16230);
   U13194 : OAI221_X1 port map( B1 => n19956, B2 => n23783, C1 => n19892, C2 =>
                           n23774, A => n16209, ZN => n16197);
   U13195 : AOI222_X1 port map( A1 => n23766, A2 => n21504, B1 => n23758, B2 =>
                           n21075, C1 => n23750, C2 => n20879, ZN => n16209);
   U13196 : OAI221_X1 port map( B1 => n19908, B2 => n23783, C1 => n19844, C2 =>
                           n23774, A => n16188, ZN => n16176);
   U13197 : AOI222_X1 port map( A1 => n23766, A2 => n21468, B1 => n23758, B2 =>
                           n21039, C1 => n23750, C2 => n20843, ZN => n16188);
   U13198 : OAI221_X1 port map( B1 => n19955, B2 => n23783, C1 => n19891, C2 =>
                           n23774, A => n16167, ZN => n16155);
   U13199 : AOI222_X1 port map( A1 => n23766, A2 => n21503, B1 => n23758, B2 =>
                           n21074, C1 => n23750, C2 => n20878, ZN => n16167);
   U13200 : OAI221_X1 port map( B1 => n19909, B2 => n23783, C1 => n19845, C2 =>
                           n23774, A => n16146, ZN => n16134);
   U13201 : AOI222_X1 port map( A1 => n23766, A2 => n21500, B1 => n23758, B2 =>
                           n21071, C1 => n23750, C2 => n20875, ZN => n16146);
   U13202 : OAI221_X1 port map( B1 => n19954, B2 => n23783, C1 => n19890, C2 =>
                           n23774, A => n16125, ZN => n16113);
   U13203 : AOI222_X1 port map( A1 => n23766, A2 => n21467, B1 => n23758, B2 =>
                           n21038, C1 => n23750, C2 => n20842, ZN => n16125);
   U13204 : OAI221_X1 port map( B1 => n19910, B2 => n23783, C1 => n19846, C2 =>
                           n23774, A => n16104, ZN => n16092);
   U13205 : AOI222_X1 port map( A1 => n23766, A2 => n21502, B1 => n23758, B2 =>
                           n21073, C1 => n23750, C2 => n20877, ZN => n16104);
   U13206 : OAI221_X1 port map( B1 => n19953, B2 => n23783, C1 => n19889, C2 =>
                           n23774, A => n16083, ZN => n16071);
   U13207 : AOI222_X1 port map( A1 => n23766, A2 => n21469, B1 => n23758, B2 =>
                           n21040, C1 => n23750, C2 => n20844, ZN => n16083);
   U13208 : OAI221_X1 port map( B1 => n19911, B2 => n23783, C1 => n19847, C2 =>
                           n23774, A => n16062, ZN => n16050);
   U13209 : AOI222_X1 port map( A1 => n23766, A2 => n21494, B1 => n23758, B2 =>
                           n21065, C1 => n23750, C2 => n20869, ZN => n16062);
   U13210 : OAI221_X1 port map( B1 => n19952, B2 => n23784, C1 => n19888, C2 =>
                           n23775, A => n16041, ZN => n16029);
   U13211 : AOI222_X1 port map( A1 => n23767, A2 => n21518, B1 => n23759, B2 =>
                           n21089, C1 => n23751, C2 => n20893, ZN => n16041);
   U13212 : OAI221_X1 port map( B1 => n19912, B2 => n23784, C1 => n19848, C2 =>
                           n23775, A => n16020, ZN => n16008);
   U13213 : AOI222_X1 port map( A1 => n23767, A2 => n21465, B1 => n23759, B2 =>
                           n21036, C1 => n23751, C2 => n20840, ZN => n16020);
   U13214 : OAI221_X1 port map( B1 => n19951, B2 => n23784, C1 => n19887, C2 =>
                           n23775, A => n15999, ZN => n15987);
   U13215 : AOI222_X1 port map( A1 => n23767, A2 => n21484, B1 => n23759, B2 =>
                           n21055, C1 => n23751, C2 => n20859, ZN => n15999);
   U13216 : OAI221_X1 port map( B1 => n19913, B2 => n23784, C1 => n19849, C2 =>
                           n23775, A => n15978, ZN => n15966);
   U13217 : AOI222_X1 port map( A1 => n23767, A2 => n21522, B1 => n23759, B2 =>
                           n21093, C1 => n23751, C2 => n20897, ZN => n15978);
   U13218 : OAI221_X1 port map( B1 => n19950, B2 => n23784, C1 => n19886, C2 =>
                           n23775, A => n15957, ZN => n15945);
   U13219 : AOI222_X1 port map( A1 => n23767, A2 => n21521, B1 => n23759, B2 =>
                           n21092, C1 => n23751, C2 => n20896, ZN => n15957);
   U13220 : OAI221_X1 port map( B1 => n19914, B2 => n23784, C1 => n19850, C2 =>
                           n23775, A => n15936, ZN => n15924);
   U13221 : AOI222_X1 port map( A1 => n23767, A2 => n21462, B1 => n23759, B2 =>
                           n21033, C1 => n23751, C2 => n20837, ZN => n15936);
   U13222 : OAI221_X1 port map( B1 => n19949, B2 => n23784, C1 => n19885, C2 =>
                           n23775, A => n15915, ZN => n15903);
   U13223 : AOI222_X1 port map( A1 => n23767, A2 => n21495, B1 => n23759, B2 =>
                           n21066, C1 => n23751, C2 => n20870, ZN => n15915);
   U13224 : OAI221_X1 port map( B1 => n19915, B2 => n23784, C1 => n19851, C2 =>
                           n23775, A => n15894, ZN => n15882);
   U13225 : AOI222_X1 port map( A1 => n23767, A2 => n21464, B1 => n23759, B2 =>
                           n21035, C1 => n23751, C2 => n20839, ZN => n15894);
   U13226 : OAI221_X1 port map( B1 => n19948, B2 => n23784, C1 => n19884, C2 =>
                           n23775, A => n15873, ZN => n15861);
   U13227 : AOI222_X1 port map( A1 => n23767, A2 => n21520, B1 => n23759, B2 =>
                           n21091, C1 => n23751, C2 => n20895, ZN => n15873);
   U13228 : OAI221_X1 port map( B1 => n19916, B2 => n23784, C1 => n19852, C2 =>
                           n23775, A => n15852, ZN => n15840);
   U13229 : AOI222_X1 port map( A1 => n23767, A2 => n21483, B1 => n23759, B2 =>
                           n21054, C1 => n23751, C2 => n20858, ZN => n15852);
   U13230 : OAI221_X1 port map( B1 => n19947, B2 => n23784, C1 => n19883, C2 =>
                           n23775, A => n15831, ZN => n15819);
   U13231 : AOI222_X1 port map( A1 => n23767, A2 => n21478, B1 => n23759, B2 =>
                           n21049, C1 => n23751, C2 => n20853, ZN => n15831);
   U13232 : OAI221_X1 port map( B1 => n19917, B2 => n23784, C1 => n19853, C2 =>
                           n23775, A => n15810, ZN => n15798);
   U13233 : AOI222_X1 port map( A1 => n23767, A2 => n21482, B1 => n23759, B2 =>
                           n21053, C1 => n23751, C2 => n20857, ZN => n15810);
   U13234 : OAI221_X1 port map( B1 => n19946, B2 => n23785, C1 => n19882, C2 =>
                           n23776, A => n15789, ZN => n15777);
   U13235 : AOI222_X1 port map( A1 => n23768, A2 => n21507, B1 => n23760, B2 =>
                           n21078, C1 => n23752, C2 => n20882, ZN => n15789);
   U13236 : OAI221_X1 port map( B1 => n19918, B2 => n23785, C1 => n19854, C2 =>
                           n23776, A => n15768, ZN => n15756);
   U13237 : AOI222_X1 port map( A1 => n23768, A2 => n21491, B1 => n23760, B2 =>
                           n21062, C1 => n23752, C2 => n20866, ZN => n15768);
   U13238 : OAI221_X1 port map( B1 => n19945, B2 => n23785, C1 => n19881, C2 =>
                           n23776, A => n15747, ZN => n15735);
   U13239 : AOI222_X1 port map( A1 => n23768, A2 => n21474, B1 => n23760, B2 =>
                           n21045, C1 => n23752, C2 => n20849, ZN => n15747);
   U13240 : OAI221_X1 port map( B1 => n19919, B2 => n23785, C1 => n19855, C2 =>
                           n23776, A => n15726, ZN => n15714);
   U13241 : AOI222_X1 port map( A1 => n23768, A2 => n21511, B1 => n23760, B2 =>
                           n21082, C1 => n23752, C2 => n20886, ZN => n15726);
   U13242 : OAI221_X1 port map( B1 => n19944, B2 => n23785, C1 => n19880, C2 =>
                           n23776, A => n15705, ZN => n15693);
   U13243 : AOI222_X1 port map( A1 => n23768, A2 => n21472, B1 => n23760, B2 =>
                           n21043, C1 => n23752, C2 => n20847, ZN => n15705);
   U13244 : OAI221_X1 port map( B1 => n19920, B2 => n23785, C1 => n19856, C2 =>
                           n23776, A => n15684, ZN => n15672);
   U13245 : AOI222_X1 port map( A1 => n23768, A2 => n21481, B1 => n23760, B2 =>
                           n21052, C1 => n23752, C2 => n20856, ZN => n15684);
   U13246 : OAI221_X1 port map( B1 => n19943, B2 => n23785, C1 => n19879, C2 =>
                           n23776, A => n15663, ZN => n15651);
   U13247 : AOI222_X1 port map( A1 => n23768, A2 => n21517, B1 => n23760, B2 =>
                           n21088, C1 => n23752, C2 => n20892, ZN => n15663);
   U13248 : OAI221_X1 port map( B1 => n19921, B2 => n23785, C1 => n19857, C2 =>
                           n23776, A => n15642, ZN => n15630);
   U13249 : AOI222_X1 port map( A1 => n23768, A2 => n21510, B1 => n23760, B2 =>
                           n21081, C1 => n23752, C2 => n20885, ZN => n15642);
   U13250 : OAI221_X1 port map( B1 => n19942, B2 => n23785, C1 => n19878, C2 =>
                           n23776, A => n15621, ZN => n15609);
   U13251 : AOI222_X1 port map( A1 => n23768, A2 => n21488, B1 => n23760, B2 =>
                           n21059, C1 => n23752, C2 => n20863, ZN => n15621);
   U13252 : OAI221_X1 port map( B1 => n19922, B2 => n23785, C1 => n19858, C2 =>
                           n23776, A => n15600, ZN => n15588);
   U13253 : AOI222_X1 port map( A1 => n23768, A2 => n21461, B1 => n23760, B2 =>
                           n21032, C1 => n23752, C2 => n20836, ZN => n15600);
   U13254 : OAI221_X1 port map( B1 => n19941, B2 => n23785, C1 => n19877, C2 =>
                           n23776, A => n15579, ZN => n15567);
   U13255 : AOI222_X1 port map( A1 => n23768, A2 => n21476, B1 => n23760, B2 =>
                           n21047, C1 => n23752, C2 => n20851, ZN => n15579);
   U13256 : OAI221_X1 port map( B1 => n19923, B2 => n23785, C1 => n19859, C2 =>
                           n23776, A => n15558, ZN => n15546);
   U13257 : AOI222_X1 port map( A1 => n23768, A2 => n21493, B1 => n23760, B2 =>
                           n21064, C1 => n23752, C2 => n20868, ZN => n15558);
   U13258 : OAI221_X1 port map( B1 => n19940, B2 => n23786, C1 => n19876, C2 =>
                           n23777, A => n15537, ZN => n15525);
   U13259 : AOI222_X1 port map( A1 => n23769, A2 => n21487, B1 => n23761, B2 =>
                           n21058, C1 => n23753, C2 => n20862, ZN => n15537);
   U13260 : OAI221_X1 port map( B1 => n19924, B2 => n23786, C1 => n19860, C2 =>
                           n23777, A => n15516, ZN => n15504);
   U13261 : AOI222_X1 port map( A1 => n23769, A2 => n21519, B1 => n23761, B2 =>
                           n21090, C1 => n23753, C2 => n20894, ZN => n15516);
   U13262 : OAI221_X1 port map( B1 => n19939, B2 => n23786, C1 => n19875, C2 =>
                           n23777, A => n15495, ZN => n15483);
   U13263 : AOI222_X1 port map( A1 => n23769, A2 => n21486, B1 => n23761, B2 =>
                           n21057, C1 => n23753, C2 => n20861, ZN => n15495);
   U13264 : OAI221_X1 port map( B1 => n19925, B2 => n23786, C1 => n19861, C2 =>
                           n23777, A => n15474, ZN => n15462);
   U13265 : AOI222_X1 port map( A1 => n23769, A2 => n21509, B1 => n23761, B2 =>
                           n21080, C1 => n23753, C2 => n20884, ZN => n15474);
   U13266 : OAI221_X1 port map( B1 => n19938, B2 => n23786, C1 => n19874, C2 =>
                           n23777, A => n15453, ZN => n15441);
   U13267 : AOI222_X1 port map( A1 => n23769, A2 => n21477, B1 => n23761, B2 =>
                           n21048, C1 => n23753, C2 => n20852, ZN => n15453);
   U13268 : OAI221_X1 port map( B1 => n19926, B2 => n23786, C1 => n19862, C2 =>
                           n23777, A => n15432, ZN => n15420);
   U13269 : AOI222_X1 port map( A1 => n23769, A2 => n21485, B1 => n23761, B2 =>
                           n21056, C1 => n23753, C2 => n20860, ZN => n15432);
   U13270 : OAI221_X1 port map( B1 => n19937, B2 => n23786, C1 => n19873, C2 =>
                           n23777, A => n15411, ZN => n15399);
   U13271 : AOI222_X1 port map( A1 => n23769, A2 => n21492, B1 => n23761, B2 =>
                           n21063, C1 => n23753, C2 => n20867, ZN => n15411);
   U13272 : OAI221_X1 port map( B1 => n19927, B2 => n23786, C1 => n19863, C2 =>
                           n23777, A => n15390, ZN => n15378);
   U13273 : AOI222_X1 port map( A1 => n23769, A2 => n21516, B1 => n23761, B2 =>
                           n21087, C1 => n23753, C2 => n20891, ZN => n15390);
   U13274 : OAI221_X1 port map( B1 => n19936, B2 => n23786, C1 => n19872, C2 =>
                           n23777, A => n15369, ZN => n15357);
   U13275 : AOI222_X1 port map( A1 => n23769, A2 => n21506, B1 => n23761, B2 =>
                           n21077, C1 => n23753, C2 => n20881, ZN => n15369);
   U13276 : OAI221_X1 port map( B1 => n19928, B2 => n23786, C1 => n19864, C2 =>
                           n23777, A => n15348, ZN => n15336);
   U13277 : AOI222_X1 port map( A1 => n23769, A2 => n21508, B1 => n23761, B2 =>
                           n21079, C1 => n23753, C2 => n20883, ZN => n15348);
   U13278 : OAI221_X1 port map( B1 => n19935, B2 => n23786, C1 => n19871, C2 =>
                           n23777, A => n15327, ZN => n15315);
   U13279 : AOI222_X1 port map( A1 => n23769, A2 => n21480, B1 => n23761, B2 =>
                           n21051, C1 => n23753, C2 => n20855, ZN => n15327);
   U13280 : OAI221_X1 port map( B1 => n19929, B2 => n23786, C1 => n19865, C2 =>
                           n23777, A => n15306, ZN => n15294);
   U13281 : AOI222_X1 port map( A1 => n23769, A2 => n21473, B1 => n23761, B2 =>
                           n21044, C1 => n23753, C2 => n20848, ZN => n15306);
   U13282 : MUX2_X1 port map( A => MEM_BUS_5_port, B => n15166, S => n23187, Z 
                           => n22701);
   U13283 : MUX2_X1 port map( A => MEM_BUS_6_port, B => n15165, S => n23187, Z 
                           => n22702);
   U13284 : MUX2_X1 port map( A => MEM_BUS_7_port, B => n15164, S => n23187, Z 
                           => n22703);
   U13285 : MUX2_X1 port map( A => MEM_BUS_8_port, B => n15163, S => n23187, Z 
                           => n22704);
   U13286 : MUX2_X1 port map( A => MEM_BUS_9_port, B => n15162, S => n23187, Z 
                           => n22705);
   U13287 : MUX2_X1 port map( A => MEM_BUS_10_port, B => n15161, S => n23187, Z
                           => n22706);
   U13288 : MUX2_X1 port map( A => MEM_BUS_11_port, B => n15160, S => n23187, Z
                           => n22707);
   U13289 : MUX2_X1 port map( A => MEM_BUS_12_port, B => n15159, S => n23188, Z
                           => n22708);
   U13290 : MUX2_X1 port map( A => MEM_BUS_13_port, B => n15158, S => n23188, Z
                           => n22709);
   U13291 : MUX2_X1 port map( A => MEM_BUS_14_port, B => n15157, S => n23188, Z
                           => n22710);
   U13292 : MUX2_X1 port map( A => MEM_BUS_15_port, B => n15156, S => n23188, Z
                           => n22711);
   U13293 : MUX2_X1 port map( A => MEM_BUS_16_port, B => n15155, S => n23188, Z
                           => n22712);
   U13294 : MUX2_X1 port map( A => MEM_BUS_17_port, B => n15154, S => n23188, Z
                           => n22713);
   U13295 : MUX2_X1 port map( A => MEM_BUS_18_port, B => n15153, S => n23188, Z
                           => n22714);
   U13296 : MUX2_X1 port map( A => MEM_BUS_19_port, B => n15152, S => n23188, Z
                           => n22715);
   U13297 : MUX2_X1 port map( A => MEM_BUS_20_port, B => n15151, S => n23188, Z
                           => n22716);
   U13298 : MUX2_X1 port map( A => MEM_BUS_21_port, B => n15150, S => n23188, Z
                           => n22717);
   U13299 : MUX2_X1 port map( A => MEM_BUS_22_port, B => n15149, S => n23188, Z
                           => n22718);
   U13300 : MUX2_X1 port map( A => MEM_BUS_23_port, B => n15148, S => n23188, Z
                           => n22719);
   U13301 : MUX2_X1 port map( A => MEM_BUS_24_port, B => n15147, S => n23189, Z
                           => n22720);
   U13302 : MUX2_X1 port map( A => MEM_BUS_25_port, B => n15146, S => n23189, Z
                           => n22721);
   U13303 : MUX2_X1 port map( A => MEM_BUS_26_port, B => n15145, S => n23189, Z
                           => n22722);
   U13304 : MUX2_X1 port map( A => MEM_BUS_27_port, B => n15144, S => n23189, Z
                           => n22723);
   U13305 : MUX2_X1 port map( A => MEM_BUS_28_port, B => n15143, S => n23189, Z
                           => n22724);
   U13306 : MUX2_X1 port map( A => MEM_BUS_29_port, B => n15142, S => n23189, Z
                           => n22725);
   U13307 : MUX2_X1 port map( A => MEM_BUS_30_port, B => n15141, S => n23189, Z
                           => n22726);
   U13308 : MUX2_X1 port map( A => MEM_BUS_31_port, B => n15140, S => n23189, Z
                           => n22727);
   U13309 : MUX2_X1 port map( A => MEM_BUS_32_port, B => n15139, S => n23189, Z
                           => n22728);
   U13310 : MUX2_X1 port map( A => MEM_BUS_33_port, B => n15138, S => n23189, Z
                           => n22729);
   U13311 : MUX2_X1 port map( A => MEM_BUS_34_port, B => n15137, S => n23189, Z
                           => n22730);
   U13312 : MUX2_X1 port map( A => MEM_BUS_35_port, B => n15136, S => n23189, Z
                           => n22731);
   U13313 : MUX2_X1 port map( A => MEM_BUS_36_port, B => n15135, S => n23190, Z
                           => n22732);
   U13314 : MUX2_X1 port map( A => MEM_BUS_37_port, B => n15134, S => n23190, Z
                           => n22733);
   U13315 : MUX2_X1 port map( A => MEM_BUS_38_port, B => n15133, S => n23190, Z
                           => n22734);
   U13316 : MUX2_X1 port map( A => MEM_BUS_39_port, B => n15132, S => n23190, Z
                           => n22735);
   U13317 : MUX2_X1 port map( A => MEM_BUS_40_port, B => n15131, S => n23190, Z
                           => n22736);
   U13318 : MUX2_X1 port map( A => MEM_BUS_41_port, B => n15130, S => n23190, Z
                           => n22737);
   U13319 : MUX2_X1 port map( A => MEM_BUS_42_port, B => n15129, S => n23190, Z
                           => n22738);
   U13320 : MUX2_X1 port map( A => MEM_BUS_43_port, B => n15128, S => n23190, Z
                           => n22739);
   U13321 : MUX2_X1 port map( A => MEM_BUS_44_port, B => n15127, S => n23190, Z
                           => n22740);
   U13322 : MUX2_X1 port map( A => MEM_BUS_45_port, B => n15126, S => n23190, Z
                           => n22741);
   U13323 : MUX2_X1 port map( A => MEM_BUS_46_port, B => n15125, S => n23190, Z
                           => n22742);
   U13324 : MUX2_X1 port map( A => MEM_BUS_47_port, B => n15124, S => n23190, Z
                           => n22743);
   U13325 : MUX2_X1 port map( A => MEM_BUS_48_port, B => n15123, S => n23191, Z
                           => n22744);
   U13326 : MUX2_X1 port map( A => MEM_BUS_49_port, B => n15122, S => n23191, Z
                           => n22745);
   U13327 : MUX2_X1 port map( A => MEM_BUS_50_port, B => n15121, S => n23191, Z
                           => n22746);
   U13328 : MUX2_X1 port map( A => MEM_BUS_51_port, B => n15120, S => n23191, Z
                           => n22747);
   U13329 : MUX2_X1 port map( A => MEM_BUS_52_port, B => n15119, S => n23191, Z
                           => n22748);
   U13330 : MUX2_X1 port map( A => MEM_BUS_53_port, B => n15118, S => n23191, Z
                           => n22749);
   U13331 : MUX2_X1 port map( A => MEM_BUS_54_port, B => n15117, S => n23191, Z
                           => n22750);
   U13332 : MUX2_X1 port map( A => MEM_BUS_55_port, B => n15116, S => n23191, Z
                           => n22751);
   U13333 : MUX2_X1 port map( A => MEM_BUS_56_port, B => n15115, S => n23191, Z
                           => n22752);
   U13334 : MUX2_X1 port map( A => MEM_BUS_57_port, B => n15114, S => n23191, Z
                           => n22753);
   U13335 : MUX2_X1 port map( A => MEM_BUS_58_port, B => n15113, S => n23191, Z
                           => n22754);
   U13336 : MUX2_X1 port map( A => MEM_BUS_59_port, B => n15112, S => n23191, Z
                           => n22755);
   U13337 : MUX2_X1 port map( A => MEM_BUS_60_port, B => n15111, S => n23192, Z
                           => n22756);
   U13338 : MUX2_X1 port map( A => MEM_BUS_61_port, B => n15110, S => n23192, Z
                           => n22757);
   U13339 : MUX2_X1 port map( A => MEM_BUS_62_port, B => n15109, S => n23192, Z
                           => n22758);
   U13340 : MUX2_X1 port map( A => MEM_BUS_63_port, B => n15108, S => n23192, Z
                           => n22759);
   U13341 : MUX2_X1 port map( A => MEM_BUS_0_port, B => n15107, S => n23187, Z 
                           => n22760);
   U13342 : NOR4_X1 port map( A1 => n15273, A2 => n15274, A3 => n15275, A4 => 
                           n15276, ZN => n15272);
   U13343 : AOI21_X1 port map( B1 => n15281, B2 => n15282, A => n23813, ZN => 
                           n15275);
   U13344 : AOI21_X1 port map( B1 => n15277, B2 => n15278, A => n23887, ZN => 
                           n15276);
   U13345 : OAI22_X1 port map( A1 => n19742, A2 => n23804, B1 => n19806, B2 => 
                           n23796, ZN => n15274);
   U13346 : NOR4_X1 port map( A1 => n15252, A2 => n15253, A3 => n15254, A4 => 
                           n15255, ZN => n15251);
   U13347 : AOI21_X1 port map( B1 => n15260, B2 => n15261, A => n23813, ZN => 
                           n15254);
   U13348 : AOI21_X1 port map( B1 => n15256, B2 => n15257, A => n23887, ZN => 
                           n15255);
   U13349 : OAI22_X1 port map( A1 => n19738, A2 => n23804, B1 => n19802, B2 => 
                           n23796, ZN => n15253);
   U13350 : NOR4_X1 port map( A1 => n15231, A2 => n15232, A3 => n15233, A4 => 
                           n15234, ZN => n15230);
   U13351 : AOI21_X1 port map( B1 => n15239, B2 => n15240, A => n23813, ZN => 
                           n15233);
   U13352 : AOI21_X1 port map( B1 => n15235, B2 => n15236, A => n23887, ZN => 
                           n15234);
   U13353 : OAI22_X1 port map( A1 => n19741, A2 => n23804, B1 => n19805, B2 => 
                           n23796, ZN => n15232);
   U13354 : NOR4_X1 port map( A1 => n15188, A2 => n15189, A3 => n15190, A4 => 
                           n15191, ZN => n15187);
   U13355 : AOI21_X1 port map( B1 => n15201, B2 => n15202, A => n23813, ZN => 
                           n15190);
   U13356 : AOI21_X1 port map( B1 => n15192, B2 => n15193, A => n23887, ZN => 
                           n15191);
   U13357 : OAI22_X1 port map( A1 => n19739, A2 => n23804, B1 => n19803, B2 => 
                           n23796, ZN => n15189);
   U13358 : OAI221_X1 port map( B1 => n19934, B2 => n23787, C1 => n19870, C2 =>
                           n23778, A => n15285, ZN => n15273);
   U13359 : AOI222_X1 port map( A1 => n23770, A2 => n21479, B1 => n23762, B2 =>
                           n21050, C1 => n23754, C2 => n20854, ZN => n15285);
   U13360 : OAI221_X1 port map( B1 => n19930, B2 => n23787, C1 => n19866, C2 =>
                           n23778, A => n15264, ZN => n15252);
   U13361 : AOI222_X1 port map( A1 => n23770, A2 => n21475, B1 => n23762, B2 =>
                           n21046, C1 => n23754, C2 => n20850, ZN => n15264);
   U13362 : OAI221_X1 port map( B1 => n19933, B2 => n23787, C1 => n19869, C2 =>
                           n23778, A => n15243, ZN => n15231);
   U13363 : AOI222_X1 port map( A1 => n23770, A2 => n21490, B1 => n23762, B2 =>
                           n21061, C1 => n23754, C2 => n20865, ZN => n15243);
   U13364 : OAI221_X1 port map( B1 => n19931, B2 => n23787, C1 => n19867, C2 =>
                           n23778, A => n15210, ZN => n15188);
   U13365 : AOI222_X1 port map( A1 => n23770, A2 => n21460, B1 => n23762, B2 =>
                           n21031, C1 => n23754, C2 => n20835, ZN => n15210);
   U13366 : MUX2_X1 port map( A => MEM_BUS_1_port, B => n15170, S => n23187, Z 
                           => n22761);
   U13367 : MUX2_X1 port map( A => MEM_BUS_2_port, B => n15169, S => n23187, Z 
                           => n22762);
   U13368 : MUX2_X1 port map( A => MEM_BUS_3_port, B => n15168, S => n23187, Z 
                           => n22763);
   U13369 : MUX2_X1 port map( A => MEM_BUS_4_port, B => n15167, S => n23187, Z 
                           => n22764);
   U13370 : OAI211_X1 port map( C1 => n3078, C2 => n23943, A => n16526, B => 
                           n16527, ZN => n5450);
   U13371 : AOI221_X1 port map( B1 => n23935, B2 => n22226, C1 => n23926, C2 =>
                           n20962, A => n16528, ZN => n16527);
   U13372 : AOI22_X1 port map( A1 => n23899, A2 => n21842, B1 => n23890, B2 => 
                           n15107, ZN => n16526);
   U13373 : OAI211_X1 port map( C1 => n3079, C2 => n23943, A => n16505, B => 
                           n16506, ZN => n5451);
   U13374 : AOI221_X1 port map( B1 => n23935, B2 => n22229, C1 => n23926, C2 =>
                           n20954, A => n16507, ZN => n16506);
   U13375 : AOI22_X1 port map( A1 => n23899, A2 => n21750, B1 => n23890, B2 => 
                           n15108, ZN => n16505);
   U13376 : OAI211_X1 port map( C1 => n3080, C2 => n23943, A => n16484, B => 
                           n16485, ZN => n5452);
   U13377 : AOI221_X1 port map( B1 => n23935, B2 => n22289, C1 => n23926, C2 =>
                           n20931, A => n16486, ZN => n16485);
   U13378 : AOI22_X1 port map( A1 => n23899, A2 => n21727, B1 => n23890, B2 => 
                           n15109, ZN => n16484);
   U13379 : OAI211_X1 port map( C1 => n3081, C2 => n23943, A => n16463, B => 
                           n16464, ZN => n5453);
   U13380 : AOI221_X1 port map( B1 => n23935, B2 => n22230, C1 => n23926, C2 =>
                           n20953, A => n16465, ZN => n16464);
   U13381 : AOI22_X1 port map( A1 => n23899, A2 => n21749, B1 => n23890, B2 => 
                           n15110, ZN => n16463);
   U13382 : OAI211_X1 port map( C1 => n3082, C2 => n23943, A => n16442, B => 
                           n16443, ZN => n5454);
   U13383 : AOI221_X1 port map( B1 => n23935, B2 => n22288, C1 => n23926, C2 =>
                           n20952, A => n16444, ZN => n16443);
   U13384 : AOI22_X1 port map( A1 => n23899, A2 => n21748, B1 => n23890, B2 => 
                           n15111, ZN => n16442);
   U13385 : OAI211_X1 port map( C1 => n3083, C2 => n23943, A => n16421, B => 
                           n16422, ZN => n5455);
   U13386 : AOI221_X1 port map( B1 => n23935, B2 => n22231, C1 => n23926, C2 =>
                           n20913, A => n16423, ZN => n16422);
   U13387 : AOI22_X1 port map( A1 => n23899, A2 => n21709, B1 => n23890, B2 => 
                           n15112, ZN => n16421);
   U13388 : OAI211_X1 port map( C1 => n3084, C2 => n23943, A => n16400, B => 
                           n16401, ZN => n5456);
   U13389 : AOI221_X1 port map( B1 => n23935, B2 => n22287, C1 => n23926, C2 =>
                           n20951, A => n16402, ZN => n16401);
   U13390 : AOI22_X1 port map( A1 => n23899, A2 => n21747, B1 => n23890, B2 => 
                           n15113, ZN => n16400);
   U13391 : OAI211_X1 port map( C1 => n3085, C2 => n23943, A => n16379, B => 
                           n16380, ZN => n5457);
   U13392 : AOI221_X1 port map( B1 => n23935, B2 => n22232, C1 => n23926, C2 =>
                           n20950, A => n16381, ZN => n16380);
   U13393 : AOI22_X1 port map( A1 => n23899, A2 => n21746, B1 => n23890, B2 => 
                           n15114, ZN => n16379);
   U13394 : OAI211_X1 port map( C1 => n3086, C2 => n23943, A => n16358, B => 
                           n16359, ZN => n5458);
   U13395 : AOI221_X1 port map( B1 => n23935, B2 => n22286, C1 => n23926, C2 =>
                           n20912, A => n16360, ZN => n16359);
   U13396 : AOI22_X1 port map( A1 => n23899, A2 => n21708, B1 => n23890, B2 => 
                           n15115, ZN => n16358);
   U13397 : OAI211_X1 port map( C1 => n3087, C2 => n23943, A => n16337, B => 
                           n16338, ZN => n5459);
   U13398 : AOI221_X1 port map( B1 => n23935, B2 => n22233, C1 => n23926, C2 =>
                           n20949, A => n16339, ZN => n16338);
   U13399 : AOI22_X1 port map( A1 => n23899, A2 => n21745, B1 => n23890, B2 => 
                           n15116, ZN => n16337);
   U13400 : OAI211_X1 port map( C1 => n3088, C2 => n23943, A => n16316, B => 
                           n16317, ZN => n5460);
   U13401 : AOI221_X1 port map( B1 => n23935, B2 => n22285, C1 => n23926, C2 =>
                           n20948, A => n16318, ZN => n16317);
   U13402 : AOI22_X1 port map( A1 => n23899, A2 => n21744, B1 => n23890, B2 => 
                           n15117, ZN => n16316);
   U13403 : OAI211_X1 port map( C1 => n3089, C2 => n23943, A => n16295, B => 
                           n16296, ZN => n5461);
   U13404 : AOI221_X1 port map( B1 => n23935, B2 => n22234, C1 => n23926, C2 =>
                           n20911, A => n16297, ZN => n16296);
   U13405 : AOI22_X1 port map( A1 => n23899, A2 => n21707, B1 => n23890, B2 => 
                           n15118, ZN => n16295);
   U13406 : OAI211_X1 port map( C1 => n3090, C2 => n23944, A => n16274, B => 
                           n16275, ZN => n5462);
   U13407 : AOI221_X1 port map( B1 => n23936, B2 => n22284, C1 => n23927, C2 =>
                           n20947, A => n16276, ZN => n16275);
   U13408 : AOI22_X1 port map( A1 => n23900, A2 => n21743, B1 => n23891, B2 => 
                           n15119, ZN => n16274);
   U13409 : OAI211_X1 port map( C1 => n3091, C2 => n23944, A => n16253, B => 
                           n16254, ZN => n5463);
   U13410 : AOI221_X1 port map( B1 => n23936, B2 => n22227, C1 => n23927, C2 =>
                           n20946, A => n16255, ZN => n16254);
   U13411 : AOI22_X1 port map( A1 => n23900, A2 => n21742, B1 => n23891, B2 => 
                           n15120, ZN => n16253);
   U13412 : OAI211_X1 port map( C1 => n3092, C2 => n23944, A => n16232, B => 
                           n16233, ZN => n5464);
   U13413 : AOI221_X1 port map( B1 => n23936, B2 => n22283, C1 => n23927, C2 =>
                           n20910, A => n16234, ZN => n16233);
   U13414 : AOI22_X1 port map( A1 => n23900, A2 => n21706, B1 => n23891, B2 => 
                           n15121, ZN => n16232);
   U13415 : OAI211_X1 port map( C1 => n3093, C2 => n23944, A => n16211, B => 
                           n16212, ZN => n5465);
   U13416 : AOI221_X1 port map( B1 => n23936, B2 => n22235, C1 => n23927, C2 =>
                           n20930, A => n16213, ZN => n16212);
   U13417 : AOI22_X1 port map( A1 => n23900, A2 => n21726, B1 => n23891, B2 => 
                           n15122, ZN => n16211);
   U13418 : OAI211_X1 port map( C1 => n3094, C2 => n23944, A => n16190, B => 
                           n16191, ZN => n5466);
   U13419 : AOI221_X1 port map( B1 => n23936, B2 => n22282, C1 => n23927, C2 =>
                           n20945, A => n16192, ZN => n16191);
   U13420 : AOI22_X1 port map( A1 => n23900, A2 => n21741, B1 => n23891, B2 => 
                           n15123, ZN => n16190);
   U13421 : OAI211_X1 port map( C1 => n3095, C2 => n23944, A => n16169, B => 
                           n16170, ZN => n5467);
   U13422 : AOI221_X1 port map( B1 => n23936, B2 => n22236, C1 => n23927, C2 =>
                           n20909, A => n16171, ZN => n16170);
   U13423 : AOI22_X1 port map( A1 => n23900, A2 => n21705, B1 => n23891, B2 => 
                           n15124, ZN => n16169);
   U13424 : OAI211_X1 port map( C1 => n3096, C2 => n23944, A => n16148, B => 
                           n16149, ZN => n5468);
   U13425 : AOI221_X1 port map( B1 => n23936, B2 => n22281, C1 => n23927, C2 =>
                           n20944, A => n16150, ZN => n16149);
   U13426 : AOI22_X1 port map( A1 => n23900, A2 => n21740, B1 => n23891, B2 => 
                           n15125, ZN => n16148);
   U13427 : OAI211_X1 port map( C1 => n3097, C2 => n23944, A => n16127, B => 
                           n16128, ZN => n5469);
   U13428 : AOI221_X1 port map( B1 => n23936, B2 => n22237, C1 => n23927, C2 =>
                           n20943, A => n16129, ZN => n16128);
   U13429 : AOI22_X1 port map( A1 => n23900, A2 => n21739, B1 => n23891, B2 => 
                           n15126, ZN => n16127);
   U13430 : OAI211_X1 port map( C1 => n3098, C2 => n23944, A => n16106, B => 
                           n16107, ZN => n5470);
   U13431 : AOI221_X1 port map( B1 => n23936, B2 => n22280, C1 => n23927, C2 =>
                           n20908, A => n16108, ZN => n16107);
   U13432 : AOI22_X1 port map( A1 => n23900, A2 => n21704, B1 => n23891, B2 => 
                           n15127, ZN => n16106);
   U13433 : OAI211_X1 port map( C1 => n3099, C2 => n23944, A => n16085, B => 
                           n16086, ZN => n5471);
   U13434 : AOI221_X1 port map( B1 => n23936, B2 => n22238, C1 => n23927, C2 =>
                           n20942, A => n16087, ZN => n16086);
   U13435 : AOI22_X1 port map( A1 => n23900, A2 => n21738, B1 => n23891, B2 => 
                           n15128, ZN => n16085);
   U13436 : OAI211_X1 port map( C1 => n3100, C2 => n23944, A => n16064, B => 
                           n16065, ZN => n5472);
   U13437 : AOI221_X1 port map( B1 => n23936, B2 => n22260, C1 => n23927, C2 =>
                           n20907, A => n16066, ZN => n16065);
   U13438 : AOI22_X1 port map( A1 => n23900, A2 => n21703, B1 => n23891, B2 => 
                           n15129, ZN => n16064);
   U13439 : OAI211_X1 port map( C1 => n3101, C2 => n23944, A => n16043, B => 
                           n16044, ZN => n5473);
   U13440 : AOI221_X1 port map( B1 => n23936, B2 => n22239, C1 => n23927, C2 =>
                           n20941, A => n16045, ZN => n16044);
   U13441 : AOI22_X1 port map( A1 => n23900, A2 => n21737, B1 => n23891, B2 => 
                           n15130, ZN => n16043);
   U13442 : OAI211_X1 port map( C1 => n3102, C2 => n23943, A => n16022, B => 
                           n16023, ZN => n5474);
   U13443 : AOI221_X1 port map( B1 => n23937, B2 => n22279, C1 => n23928, C2 =>
                           n20958, A => n16024, ZN => n16023);
   U13444 : AOI22_X1 port map( A1 => n23901, A2 => n21836, B1 => n23892, B2 => 
                           n15131, ZN => n16022);
   U13445 : OAI211_X1 port map( C1 => n3103, C2 => n23944, A => n16001, B => 
                           n16002, ZN => n5475);
   U13446 : AOI221_X1 port map( B1 => n23937, B2 => n22240, C1 => n23928, C2 =>
                           n20906, A => n16003, ZN => n16002);
   U13447 : AOI22_X1 port map( A1 => n23901, A2 => n21702, B1 => n23892, B2 => 
                           n15132, ZN => n16001);
   U13448 : OAI211_X1 port map( C1 => n3104, C2 => n23943, A => n15980, B => 
                           n15981, ZN => n5476);
   U13449 : AOI221_X1 port map( B1 => n23937, B2 => n22278, C1 => n23928, C2 =>
                           n20929, A => n15982, ZN => n15981);
   U13450 : AOI22_X1 port map( A1 => n23901, A2 => n21725, B1 => n23892, B2 => 
                           n15133, ZN => n15980);
   U13451 : OAI211_X1 port map( C1 => n3105, C2 => n23944, A => n15959, B => 
                           n15960, ZN => n5477);
   U13452 : AOI221_X1 port map( B1 => n23937, B2 => n22241, C1 => n23928, C2 =>
                           n20961, A => n15961, ZN => n15960);
   U13453 : AOI22_X1 port map( A1 => n23901, A2 => n21839, B1 => n23892, B2 => 
                           n15134, ZN => n15959);
   U13454 : OAI211_X1 port map( C1 => n3106, C2 => n23945, A => n15938, B => 
                           n15939, ZN => n5478);
   U13455 : AOI221_X1 port map( B1 => n23937, B2 => n22277, C1 => n23928, C2 =>
                           n20960, A => n15940, ZN => n15939);
   U13456 : AOI22_X1 port map( A1 => n23901, A2 => n21838, B1 => n23892, B2 => 
                           n15135, ZN => n15938);
   U13457 : OAI211_X1 port map( C1 => n3107, C2 => n23945, A => n15917, B => 
                           n15918, ZN => n5479);
   U13458 : AOI221_X1 port map( B1 => n23937, B2 => n22242, C1 => n23928, C2 =>
                           n20905, A => n15919, ZN => n15918);
   U13459 : AOI22_X1 port map( A1 => n23901, A2 => n21701, B1 => n23892, B2 => 
                           n15136, ZN => n15917);
   U13460 : OAI211_X1 port map( C1 => n3108, C2 => n23945, A => n15896, B => 
                           n15897, ZN => n5480);
   U13461 : AOI221_X1 port map( B1 => n23937, B2 => n22276, C1 => n23928, C2 =>
                           n20940, A => n15898, ZN => n15897);
   U13462 : AOI22_X1 port map( A1 => n23901, A2 => n21736, B1 => n23892, B2 => 
                           n15137, ZN => n15896);
   U13463 : OAI211_X1 port map( C1 => n3109, C2 => n23945, A => n15875, B => 
                           n15876, ZN => n5481);
   U13464 : AOI221_X1 port map( B1 => n23937, B2 => n22243, C1 => n23928, C2 =>
                           n20904, A => n15877, ZN => n15876);
   U13465 : AOI22_X1 port map( A1 => n23901, A2 => n21700, B1 => n23892, B2 => 
                           n15138, ZN => n15875);
   U13466 : OAI211_X1 port map( C1 => n3110, C2 => n23945, A => n15854, B => 
                           n15855, ZN => n5482);
   U13467 : AOI221_X1 port map( B1 => n23937, B2 => n22275, C1 => n23928, C2 =>
                           n20959, A => n15856, ZN => n15855);
   U13468 : AOI22_X1 port map( A1 => n23901, A2 => n21837, B1 => n23892, B2 => 
                           n15139, ZN => n15854);
   U13469 : OAI211_X1 port map( C1 => n3111, C2 => n23945, A => n15833, B => 
                           n15834, ZN => n5483);
   U13470 : AOI221_X1 port map( B1 => n23937, B2 => n22244, C1 => n23928, C2 =>
                           n20928, A => n15835, ZN => n15834);
   U13471 : AOI22_X1 port map( A1 => n23901, A2 => n21724, B1 => n23892, B2 => 
                           n15140, ZN => n15833);
   U13472 : OAI211_X1 port map( C1 => n3112, C2 => n23945, A => n15812, B => 
                           n15813, ZN => n5484);
   U13473 : AOI221_X1 port map( B1 => n23937, B2 => n22274, C1 => n23928, C2 =>
                           n20927, A => n15814, ZN => n15813);
   U13474 : AOI22_X1 port map( A1 => n23901, A2 => n21723, B1 => n23892, B2 => 
                           n15141, ZN => n15812);
   U13475 : OAI211_X1 port map( C1 => n3113, C2 => n23945, A => n15791, B => 
                           n15792, ZN => n5485);
   U13476 : AOI221_X1 port map( B1 => n23937, B2 => n22245, C1 => n23928, C2 =>
                           n20926, A => n15793, ZN => n15792);
   U13477 : AOI22_X1 port map( A1 => n23901, A2 => n21722, B1 => n23892, B2 => 
                           n15142, ZN => n15791);
   U13478 : OAI211_X1 port map( C1 => n3114, C2 => n23943, A => n15770, B => 
                           n15771, ZN => n5486);
   U13479 : AOI221_X1 port map( B1 => n23938, B2 => n22273, C1 => n23929, C2 =>
                           n20939, A => n15772, ZN => n15771);
   U13480 : AOI22_X1 port map( A1 => n23902, A2 => n21735, B1 => n23893, B2 => 
                           n15143, ZN => n15770);
   U13481 : OAI211_X1 port map( C1 => n3115, C2 => n23944, A => n15749, B => 
                           n15750, ZN => n5487);
   U13482 : AOI221_X1 port map( B1 => n23938, B2 => n22228, C1 => n23929, C2 =>
                           n20925, A => n15751, ZN => n15750);
   U13483 : AOI22_X1 port map( A1 => n23902, A2 => n21721, B1 => n23893, B2 => 
                           n15144, ZN => n15749);
   U13484 : OAI211_X1 port map( C1 => n3116, C2 => n23944, A => n15728, B => 
                           n15729, ZN => n5488);
   U13485 : AOI221_X1 port map( B1 => n23938, B2 => n22272, C1 => n23929, C2 =>
                           n20903, A => n15730, ZN => n15729);
   U13486 : AOI22_X1 port map( A1 => n23902, A2 => n21699, B1 => n23893, B2 => 
                           n15145, ZN => n15728);
   U13487 : OAI211_X1 port map( C1 => n3117, C2 => n23943, A => n15707, B => 
                           n15708, ZN => n5489);
   U13488 : AOI221_X1 port map( B1 => n23938, B2 => n22246, C1 => n23929, C2 =>
                           n20938, A => n15709, ZN => n15708);
   U13489 : AOI22_X1 port map( A1 => n23902, A2 => n21734, B1 => n23893, B2 => 
                           n15146, ZN => n15707);
   U13490 : OAI211_X1 port map( C1 => n3118, C2 => n23944, A => n15686, B => 
                           n15687, ZN => n5490);
   U13491 : AOI221_X1 port map( B1 => n23938, B2 => n22271, C1 => n23929, C2 =>
                           n20899, A => n15688, ZN => n15687);
   U13492 : AOI22_X1 port map( A1 => n23902, A2 => n21698, B1 => n23893, B2 => 
                           n15147, ZN => n15686);
   U13493 : OAI211_X1 port map( C1 => n3119, C2 => n23943, A => n15665, B => 
                           n15666, ZN => n5491);
   U13494 : AOI221_X1 port map( B1 => n23938, B2 => n22247, C1 => n23929, C2 =>
                           n20924, A => n15667, ZN => n15666);
   U13495 : AOI22_X1 port map( A1 => n23902, A2 => n21720, B1 => n23893, B2 => 
                           n15148, ZN => n15665);
   U13496 : OAI211_X1 port map( C1 => n3120, C2 => n23943, A => n15644, B => 
                           n15645, ZN => n5492);
   U13497 : AOI221_X1 port map( B1 => n23938, B2 => n22270, C1 => n23929, C2 =>
                           n20956, A => n15646, ZN => n15645);
   U13498 : AOI22_X1 port map( A1 => n23902, A2 => n21765, B1 => n23893, B2 => 
                           n15149, ZN => n15644);
   U13499 : OAI211_X1 port map( C1 => n3121, C2 => n23944, A => n15623, B => 
                           n15624, ZN => n5493);
   U13500 : AOI221_X1 port map( B1 => n23938, B2 => n22248, C1 => n23929, C2 =>
                           n20937, A => n15625, ZN => n15624);
   U13501 : AOI22_X1 port map( A1 => n23902, A2 => n21733, B1 => n23893, B2 => 
                           n15150, ZN => n15623);
   U13502 : OAI211_X1 port map( C1 => n3122, C2 => n23944, A => n15602, B => 
                           n15603, ZN => n5494);
   U13503 : AOI221_X1 port map( B1 => n23938, B2 => n22269, C1 => n23929, C2 =>
                           n20923, A => n15604, ZN => n15603);
   U13504 : AOI22_X1 port map( A1 => n23902, A2 => n21719, B1 => n23893, B2 => 
                           n15151, ZN => n15602);
   U13505 : OAI211_X1 port map( C1 => n3123, C2 => n23943, A => n15581, B => 
                           n15582, ZN => n5495);
   U13506 : AOI221_X1 port map( B1 => n23938, B2 => n22249, C1 => n23929, C2 =>
                           n20902, A => n15583, ZN => n15582);
   U13507 : AOI22_X1 port map( A1 => n23902, A2 => n21697, B1 => n23893, B2 => 
                           n15152, ZN => n15581);
   U13508 : OAI211_X1 port map( C1 => n3124, C2 => n23944, A => n15560, B => 
                           n15561, ZN => n5496);
   U13509 : AOI221_X1 port map( B1 => n23938, B2 => n22259, C1 => n23929, C2 =>
                           n20922, A => n15562, ZN => n15561);
   U13510 : AOI22_X1 port map( A1 => n23902, A2 => n21718, B1 => n23893, B2 => 
                           n15153, ZN => n15560);
   U13511 : OAI211_X1 port map( C1 => n3125, C2 => n23943, A => n15539, B => 
                           n15540, ZN => n5497);
   U13512 : AOI221_X1 port map( B1 => n23938, B2 => n22261, C1 => n23929, C2 =>
                           n20936, A => n15541, ZN => n15540);
   U13513 : AOI22_X1 port map( A1 => n23902, A2 => n21732, B1 => n23893, B2 => 
                           n15154, ZN => n15539);
   U13514 : OAI211_X1 port map( C1 => n3126, C2 => n23943, A => n15518, B => 
                           n15519, ZN => n5498);
   U13515 : AOI221_X1 port map( B1 => n23939, B2 => n22268, C1 => n23930, C2 =>
                           n20921, A => n15520, ZN => n15519);
   U13516 : AOI22_X1 port map( A1 => n23903, A2 => n21717, B1 => n23894, B2 => 
                           n15155, ZN => n15518);
   U13517 : OAI211_X1 port map( C1 => n3127, C2 => n23943, A => n15497, B => 
                           n15498, ZN => n5499);
   U13518 : AOI221_X1 port map( B1 => n23939, B2 => n22250, C1 => n23930, C2 =>
                           n20957, A => n15499, ZN => n15498);
   U13519 : AOI22_X1 port map( A1 => n23903, A2 => n21835, B1 => n23894, B2 => 
                           n15156, ZN => n15497);
   U13520 : OAI211_X1 port map( C1 => n3128, C2 => n23944, A => n15476, B => 
                           n15477, ZN => n5500);
   U13521 : AOI221_X1 port map( B1 => n23939, B2 => n22267, C1 => n23930, C2 =>
                           n20920, A => n15478, ZN => n15477);
   U13522 : AOI22_X1 port map( A1 => n23903, A2 => n21716, B1 => n23894, B2 => 
                           n15157, ZN => n15476);
   U13523 : OAI211_X1 port map( C1 => n3129, C2 => n23944, A => n15455, B => 
                           n15456, ZN => n5501);
   U13524 : AOI221_X1 port map( B1 => n23939, B2 => n22251, C1 => n23930, C2 =>
                           n20935, A => n15457, ZN => n15456);
   U13525 : AOI22_X1 port map( A1 => n23903, A2 => n21731, B1 => n23894, B2 => 
                           n15158, ZN => n15455);
   U13526 : OAI211_X1 port map( C1 => n3130, C2 => n23944, A => n15434, B => 
                           n15435, ZN => n5502);
   U13527 : AOI221_X1 port map( B1 => n23939, B2 => n22266, C1 => n23930, C2 =>
                           n20919, A => n15436, ZN => n15435);
   U13528 : AOI22_X1 port map( A1 => n23903, A2 => n21715, B1 => n23894, B2 => 
                           n15159, ZN => n15434);
   U13529 : OAI211_X1 port map( C1 => n3131, C2 => n23943, A => n15413, B => 
                           n15414, ZN => n5503);
   U13530 : AOI221_X1 port map( B1 => n23939, B2 => n22252, C1 => n23930, C2 =>
                           n20918, A => n15415, ZN => n15414);
   U13531 : AOI22_X1 port map( A1 => n23903, A2 => n21714, B1 => n23894, B2 => 
                           n15160, ZN => n15413);
   U13532 : OAI211_X1 port map( C1 => n3132, C2 => n23944, A => n15392, B => 
                           n15393, ZN => n5504);
   U13533 : AOI221_X1 port map( B1 => n23939, B2 => n22265, C1 => n23930, C2 =>
                           n20934, A => n15394, ZN => n15393);
   U13534 : AOI22_X1 port map( A1 => n23903, A2 => n21730, B1 => n23894, B2 => 
                           n15161, ZN => n15392);
   U13535 : OAI211_X1 port map( C1 => n3133, C2 => n23943, A => n15371, B => 
                           n15372, ZN => n5505);
   U13536 : AOI221_X1 port map( B1 => n23939, B2 => n22253, C1 => n23930, C2 =>
                           n20955, A => n15373, ZN => n15372);
   U13537 : AOI22_X1 port map( A1 => n23903, A2 => n21754, B1 => n23894, B2 => 
                           n15162, ZN => n15371);
   U13538 : OAI211_X1 port map( C1 => n3134, C2 => n23943, A => n15350, B => 
                           n15351, ZN => n5506);
   U13539 : AOI221_X1 port map( B1 => n23939, B2 => n22264, C1 => n23930, C2 =>
                           n20933, A => n15352, ZN => n15351);
   U13540 : AOI22_X1 port map( A1 => n23903, A2 => n21729, B1 => n23894, B2 => 
                           n15163, ZN => n15350);
   U13541 : OAI211_X1 port map( C1 => n3135, C2 => n23943, A => n15329, B => 
                           n15330, ZN => n5507);
   U13542 : AOI221_X1 port map( B1 => n23939, B2 => n22254, C1 => n23930, C2 =>
                           n20932, A => n15331, ZN => n15330);
   U13543 : AOI22_X1 port map( A1 => n23903, A2 => n21728, B1 => n23894, B2 => 
                           n15164, ZN => n15329);
   U13544 : OAI211_X1 port map( C1 => n3136, C2 => n23944, A => n15308, B => 
                           n15309, ZN => n5508);
   U13545 : AOI221_X1 port map( B1 => n23939, B2 => n22263, C1 => n23930, C2 =>
                           n20917, A => n15310, ZN => n15309);
   U13546 : AOI22_X1 port map( A1 => n23903, A2 => n21713, B1 => n23894, B2 => 
                           n15165, ZN => n15308);
   U13547 : OAI211_X1 port map( C1 => n3137, C2 => n23944, A => n15287, B => 
                           n15288, ZN => n5509);
   U13548 : AOI221_X1 port map( B1 => n23939, B2 => n22262, C1 => n23930, C2 =>
                           n20901, A => n15289, ZN => n15288);
   U13549 : AOI22_X1 port map( A1 => n23903, A2 => n21696, B1 => n23894, B2 => 
                           n15166, ZN => n15287);
   U13550 : OAI211_X1 port map( C1 => n3138, C2 => n23945, A => n15266, B => 
                           n15267, ZN => n5510);
   U13551 : AOI221_X1 port map( B1 => n23940, B2 => n22258, C1 => n23931, C2 =>
                           n20916, A => n15268, ZN => n15267);
   U13552 : AOI22_X1 port map( A1 => n23904, A2 => n21712, B1 => n23895, B2 => 
                           n15167, ZN => n15266);
   U13553 : OAI211_X1 port map( C1 => n3139, C2 => n23945, A => n15245, B => 
                           n15246, ZN => n5511);
   U13554 : AOI221_X1 port map( B1 => n23940, B2 => n22255, C1 => n23931, C2 =>
                           n20915, A => n15247, ZN => n15246);
   U13555 : AOI22_X1 port map( A1 => n23904, A2 => n21711, B1 => n23895, B2 => 
                           n15168, ZN => n15245);
   U13556 : OAI211_X1 port map( C1 => n3140, C2 => n23945, A => n15224, B => 
                           n15225, ZN => n5512);
   U13557 : AOI221_X1 port map( B1 => n23940, B2 => n22257, C1 => n23931, C2 =>
                           n20914, A => n15226, ZN => n15225);
   U13558 : AOI22_X1 port map( A1 => n23904, A2 => n21710, B1 => n23895, B2 => 
                           n15169, ZN => n15224);
   U13559 : OAI211_X1 port map( C1 => n3141, C2 => n23945, A => n15175, B => 
                           n15176, ZN => n5513);
   U13560 : AOI221_X1 port map( B1 => n23940, B2 => n22256, C1 => n23931, C2 =>
                           n20900, A => n15179, ZN => n15176);
   U13561 : AOI22_X1 port map( A1 => n23904, A2 => n21695, B1 => n23895, B2 => 
                           n15170, ZN => n15175);
   U13562 : OAI22_X1 port map( A1 => n20188, A2 => n23723, B1 => n20252, B2 => 
                           n23714, ZN => n16554);
   U13563 : OAI22_X1 port map( A1 => n20156, A2 => n23723, B1 => n20220, B2 => 
                           n23714, ZN => n16525);
   U13564 : OAI22_X1 port map( A1 => n20219, A2 => n23723, B1 => n20283, B2 => 
                           n23714, ZN => n16504);
   U13565 : OAI22_X1 port map( A1 => n20157, A2 => n23723, B1 => n20221, B2 => 
                           n23714, ZN => n16483);
   U13566 : OAI22_X1 port map( A1 => n20218, A2 => n23723, B1 => n20282, B2 => 
                           n23714, ZN => n16462);
   U13567 : OAI22_X1 port map( A1 => n20158, A2 => n23723, B1 => n20222, B2 => 
                           n23714, ZN => n16441);
   U13568 : OAI22_X1 port map( A1 => n20217, A2 => n23723, B1 => n20281, B2 => 
                           n23714, ZN => n16420);
   U13569 : OAI22_X1 port map( A1 => n20159, A2 => n23723, B1 => n20223, B2 => 
                           n23714, ZN => n16399);
   U13570 : OAI22_X1 port map( A1 => n20216, A2 => n23723, B1 => n20280, B2 => 
                           n23714, ZN => n16378);
   U13571 : OAI22_X1 port map( A1 => n20160, A2 => n23723, B1 => n20224, B2 => 
                           n23714, ZN => n16357);
   U13572 : OAI22_X1 port map( A1 => n20215, A2 => n23723, B1 => n20279, B2 => 
                           n23714, ZN => n16336);
   U13573 : OAI22_X1 port map( A1 => n20161, A2 => n23723, B1 => n20225, B2 => 
                           n23714, ZN => n16315);
   U13574 : OAI22_X1 port map( A1 => n20214, A2 => n23724, B1 => n20278, B2 => 
                           n23715, ZN => n16294);
   U13575 : OAI22_X1 port map( A1 => n20162, A2 => n23724, B1 => n20226, B2 => 
                           n23715, ZN => n16273);
   U13576 : OAI22_X1 port map( A1 => n20213, A2 => n23724, B1 => n20277, B2 => 
                           n23715, ZN => n16252);
   U13577 : OAI22_X1 port map( A1 => n20163, A2 => n23724, B1 => n20227, B2 => 
                           n23715, ZN => n16231);
   U13578 : OAI22_X1 port map( A1 => n20212, A2 => n23724, B1 => n20276, B2 => 
                           n23715, ZN => n16210);
   U13579 : OAI22_X1 port map( A1 => n20164, A2 => n23724, B1 => n20228, B2 => 
                           n23715, ZN => n16189);
   U13580 : OAI22_X1 port map( A1 => n20211, A2 => n23724, B1 => n20275, B2 => 
                           n23715, ZN => n16168);
   U13581 : OAI22_X1 port map( A1 => n20165, A2 => n23724, B1 => n20229, B2 => 
                           n23715, ZN => n16147);
   U13582 : OAI22_X1 port map( A1 => n20210, A2 => n23724, B1 => n20274, B2 => 
                           n23715, ZN => n16126);
   U13583 : OAI22_X1 port map( A1 => n20166, A2 => n23724, B1 => n20230, B2 => 
                           n23715, ZN => n16105);
   U13584 : OAI22_X1 port map( A1 => n20209, A2 => n23724, B1 => n20273, B2 => 
                           n23715, ZN => n16084);
   U13585 : OAI22_X1 port map( A1 => n20167, A2 => n23724, B1 => n20231, B2 => 
                           n23715, ZN => n16063);
   U13586 : OAI22_X1 port map( A1 => n20208, A2 => n23725, B1 => n20272, B2 => 
                           n23716, ZN => n16042);
   U13587 : OAI22_X1 port map( A1 => n20168, A2 => n23725, B1 => n20232, B2 => 
                           n23716, ZN => n16021);
   U13588 : OAI22_X1 port map( A1 => n20207, A2 => n23725, B1 => n20271, B2 => 
                           n23716, ZN => n16000);
   U13589 : OAI22_X1 port map( A1 => n20169, A2 => n23725, B1 => n20233, B2 => 
                           n23716, ZN => n15979);
   U13590 : OAI22_X1 port map( A1 => n20206, A2 => n23725, B1 => n20270, B2 => 
                           n23716, ZN => n15958);
   U13591 : OAI22_X1 port map( A1 => n20170, A2 => n23725, B1 => n20234, B2 => 
                           n23716, ZN => n15937);
   U13592 : OAI22_X1 port map( A1 => n20205, A2 => n23725, B1 => n20269, B2 => 
                           n23716, ZN => n15916);
   U13593 : OAI22_X1 port map( A1 => n20171, A2 => n23725, B1 => n20235, B2 => 
                           n23716, ZN => n15895);
   U13594 : OAI22_X1 port map( A1 => n20204, A2 => n23725, B1 => n20268, B2 => 
                           n23716, ZN => n15874);
   U13595 : OAI22_X1 port map( A1 => n20172, A2 => n23725, B1 => n20236, B2 => 
                           n23716, ZN => n15853);
   U13596 : OAI22_X1 port map( A1 => n20203, A2 => n23725, B1 => n20267, B2 => 
                           n23716, ZN => n15832);
   U13597 : OAI22_X1 port map( A1 => n20173, A2 => n23725, B1 => n20237, B2 => 
                           n23716, ZN => n15811);
   U13598 : OAI22_X1 port map( A1 => n20202, A2 => n23726, B1 => n20266, B2 => 
                           n23717, ZN => n15790);
   U13599 : OAI22_X1 port map( A1 => n20174, A2 => n23726, B1 => n20238, B2 => 
                           n23717, ZN => n15769);
   U13600 : OAI22_X1 port map( A1 => n20201, A2 => n23726, B1 => n20265, B2 => 
                           n23717, ZN => n15748);
   U13601 : OAI22_X1 port map( A1 => n20175, A2 => n23726, B1 => n20239, B2 => 
                           n23717, ZN => n15727);
   U13602 : OAI22_X1 port map( A1 => n20200, A2 => n23726, B1 => n20264, B2 => 
                           n23717, ZN => n15706);
   U13603 : OAI22_X1 port map( A1 => n20176, A2 => n23726, B1 => n20240, B2 => 
                           n23717, ZN => n15685);
   U13604 : OAI22_X1 port map( A1 => n20199, A2 => n23726, B1 => n20263, B2 => 
                           n23717, ZN => n15664);
   U13605 : OAI22_X1 port map( A1 => n20177, A2 => n23726, B1 => n20241, B2 => 
                           n23717, ZN => n15643);
   U13606 : OAI22_X1 port map( A1 => n20198, A2 => n23726, B1 => n20262, B2 => 
                           n23717, ZN => n15622);
   U13607 : OAI22_X1 port map( A1 => n20178, A2 => n23726, B1 => n20242, B2 => 
                           n23717, ZN => n15601);
   U13608 : OAI22_X1 port map( A1 => n20197, A2 => n23726, B1 => n20261, B2 => 
                           n23717, ZN => n15580);
   U13609 : OAI22_X1 port map( A1 => n20179, A2 => n23726, B1 => n20243, B2 => 
                           n23717, ZN => n15559);
   U13610 : OAI22_X1 port map( A1 => n20196, A2 => n23727, B1 => n20260, B2 => 
                           n23718, ZN => n15538);
   U13611 : OAI22_X1 port map( A1 => n20180, A2 => n23727, B1 => n20244, B2 => 
                           n23718, ZN => n15517);
   U13612 : OAI22_X1 port map( A1 => n20195, A2 => n23727, B1 => n20259, B2 => 
                           n23718, ZN => n15496);
   U13613 : OAI22_X1 port map( A1 => n20181, A2 => n23727, B1 => n20245, B2 => 
                           n23718, ZN => n15475);
   U13614 : OAI22_X1 port map( A1 => n20194, A2 => n23727, B1 => n20258, B2 => 
                           n23718, ZN => n15454);
   U13615 : OAI22_X1 port map( A1 => n20182, A2 => n23727, B1 => n20246, B2 => 
                           n23718, ZN => n15433);
   U13616 : OAI22_X1 port map( A1 => n20193, A2 => n23727, B1 => n20257, B2 => 
                           n23718, ZN => n15412);
   U13617 : OAI22_X1 port map( A1 => n20183, A2 => n23727, B1 => n20247, B2 => 
                           n23718, ZN => n15391);
   U13618 : OAI22_X1 port map( A1 => n20192, A2 => n23727, B1 => n20256, B2 => 
                           n23718, ZN => n15370);
   U13619 : OAI22_X1 port map( A1 => n20184, A2 => n23727, B1 => n20248, B2 => 
                           n23718, ZN => n15349);
   U13620 : OAI22_X1 port map( A1 => n20191, A2 => n23727, B1 => n20255, B2 => 
                           n23718, ZN => n15328);
   U13621 : OAI22_X1 port map( A1 => n20185, A2 => n23727, B1 => n20249, B2 => 
                           n23718, ZN => n15307);
   U13622 : OAI22_X1 port map( A1 => n20190, A2 => n23728, B1 => n20254, B2 => 
                           n23719, ZN => n15286);
   U13623 : OAI22_X1 port map( A1 => n20186, A2 => n23728, B1 => n20250, B2 => 
                           n23719, ZN => n15265);
   U13624 : OAI22_X1 port map( A1 => n20189, A2 => n23728, B1 => n20253, B2 => 
                           n23719, ZN => n15244);
   U13625 : OAI22_X1 port map( A1 => n20187, A2 => n23728, B1 => n20251, B2 => 
                           n23719, ZN => n15216);
   U13626 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => n22768, ZN => n22765);
   U13627 : OAI22_X1 port map( A1 => n16635, A2 => n23522, B1 => n20638, B2 => 
                           n22821, ZN => n3460);
   U13628 : OAI22_X1 port map( A1 => n16634, A2 => n23522, B1 => n20637, B2 => 
                           n22821, ZN => n3461);
   U13629 : OAI22_X1 port map( A1 => n16633, A2 => n23522, B1 => n20636, B2 => 
                           n22821, ZN => n3462);
   U13630 : OAI22_X1 port map( A1 => n16632, A2 => n23522, B1 => n20635, B2 => 
                           n22821, ZN => n3463);
   U13631 : OAI22_X1 port map( A1 => n16631, A2 => n23522, B1 => n20634, B2 => 
                           n22821, ZN => n3464);
   U13632 : OAI22_X1 port map( A1 => n16630, A2 => n23522, B1 => n20633, B2 => 
                           n22821, ZN => n3465);
   U13633 : OAI22_X1 port map( A1 => n16629, A2 => n23522, B1 => n20632, B2 => 
                           n22821, ZN => n3466);
   U13634 : OAI22_X1 port map( A1 => n16623, A2 => n23524, B1 => n20626, B2 => 
                           n22822, ZN => n3472);
   U13635 : OAI22_X1 port map( A1 => n16622, A2 => n23523, B1 => n20625, B2 => 
                           n22822, ZN => n3473);
   U13636 : OAI22_X1 port map( A1 => n16621, A2 => n23522, B1 => n20624, B2 => 
                           n22822, ZN => n3474);
   U13637 : OAI22_X1 port map( A1 => n16620, A2 => n23524, B1 => n20623, B2 => 
                           n22822, ZN => n3475);
   U13638 : OAI22_X1 port map( A1 => n16619, A2 => n23523, B1 => n20622, B2 => 
                           n22822, ZN => n3476);
   U13639 : OAI22_X1 port map( A1 => n16618, A2 => n23522, B1 => n20621, B2 => 
                           n22822, ZN => n3477);
   U13640 : OAI22_X1 port map( A1 => n16617, A2 => n23524, B1 => n20620, B2 => 
                           n22822, ZN => n3478);
   U13641 : OAI22_X1 port map( A1 => n16611, A2 => n23522, B1 => n20614, B2 => 
                           n22823, ZN => n3484);
   U13642 : OAI22_X1 port map( A1 => n16610, A2 => n23522, B1 => n20613, B2 => 
                           n22823, ZN => n3485);
   U13643 : OAI22_X1 port map( A1 => n16609, A2 => n23524, B1 => n20612, B2 => 
                           n22823, ZN => n3486);
   U13644 : OAI22_X1 port map( A1 => n16608, A2 => n23523, B1 => n20611, B2 => 
                           n22823, ZN => n3487);
   U13645 : OAI22_X1 port map( A1 => n16607, A2 => n23522, B1 => n20610, B2 => 
                           n22823, ZN => n3488);
   U13646 : OAI22_X1 port map( A1 => n16606, A2 => n23522, B1 => n20609, B2 => 
                           n22823, ZN => n3489);
   U13647 : OAI22_X1 port map( A1 => n16605, A2 => n23524, B1 => n20608, B2 => 
                           n22823, ZN => n3490);
   U13648 : OAI22_X1 port map( A1 => n16635, A2 => n23542, B1 => n20510, B2 => 
                           n22833, ZN => n3588);
   U13649 : OAI22_X1 port map( A1 => n16634, A2 => n23542, B1 => n20509, B2 => 
                           n22833, ZN => n3589);
   U13650 : OAI22_X1 port map( A1 => n16633, A2 => n23542, B1 => n20508, B2 => 
                           n22833, ZN => n3590);
   U13651 : OAI22_X1 port map( A1 => n16632, A2 => n23542, B1 => n20507, B2 => 
                           n22833, ZN => n3591);
   U13652 : OAI22_X1 port map( A1 => n16631, A2 => n23542, B1 => n20506, B2 => 
                           n22833, ZN => n3592);
   U13653 : OAI22_X1 port map( A1 => n16630, A2 => n23542, B1 => n20505, B2 => 
                           n22833, ZN => n3593);
   U13654 : OAI22_X1 port map( A1 => n16629, A2 => n23542, B1 => n20504, B2 => 
                           n22833, ZN => n3594);
   U13655 : OAI22_X1 port map( A1 => n16623, A2 => n23544, B1 => n20498, B2 => 
                           n22834, ZN => n3600);
   U13656 : OAI22_X1 port map( A1 => n16622, A2 => n23543, B1 => n20497, B2 => 
                           n22834, ZN => n3601);
   U13657 : OAI22_X1 port map( A1 => n16621, A2 => n23542, B1 => n20496, B2 => 
                           n22834, ZN => n3602);
   U13658 : OAI22_X1 port map( A1 => n16620, A2 => n23544, B1 => n20495, B2 => 
                           n22834, ZN => n3603);
   U13659 : OAI22_X1 port map( A1 => n16619, A2 => n23543, B1 => n20494, B2 => 
                           n22834, ZN => n3604);
   U13660 : OAI22_X1 port map( A1 => n16618, A2 => n23542, B1 => n20493, B2 => 
                           n22834, ZN => n3605);
   U13661 : OAI22_X1 port map( A1 => n16617, A2 => n23544, B1 => n20492, B2 => 
                           n22834, ZN => n3606);
   U13662 : OAI22_X1 port map( A1 => n16611, A2 => n23542, B1 => n20486, B2 => 
                           n22835, ZN => n3612);
   U13663 : OAI22_X1 port map( A1 => n16610, A2 => n23542, B1 => n20485, B2 => 
                           n22835, ZN => n3613);
   U13664 : OAI22_X1 port map( A1 => n16609, A2 => n23544, B1 => n20484, B2 => 
                           n22835, ZN => n3614);
   U13665 : OAI22_X1 port map( A1 => n16608, A2 => n23543, B1 => n20483, B2 => 
                           n22835, ZN => n3615);
   U13666 : OAI22_X1 port map( A1 => n16607, A2 => n23542, B1 => n20482, B2 => 
                           n22835, ZN => n3616);
   U13667 : OAI22_X1 port map( A1 => n16606, A2 => n23542, B1 => n20481, B2 => 
                           n22835, ZN => n3617);
   U13668 : OAI22_X1 port map( A1 => n16605, A2 => n23544, B1 => n20480, B2 => 
                           n22835, ZN => n3618);
   U13669 : OAI22_X1 port map( A1 => n16635, A2 => n23562, B1 => n20382, B2 => 
                           n22845, ZN => n3716);
   U13670 : OAI22_X1 port map( A1 => n16634, A2 => n23562, B1 => n20381, B2 => 
                           n22845, ZN => n3717);
   U13671 : OAI22_X1 port map( A1 => n16633, A2 => n23562, B1 => n20380, B2 => 
                           n22845, ZN => n3718);
   U13672 : OAI22_X1 port map( A1 => n16632, A2 => n23562, B1 => n20379, B2 => 
                           n22845, ZN => n3719);
   U13673 : OAI22_X1 port map( A1 => n16631, A2 => n23562, B1 => n20378, B2 => 
                           n22845, ZN => n3720);
   U13674 : OAI22_X1 port map( A1 => n16630, A2 => n23562, B1 => n20377, B2 => 
                           n22845, ZN => n3721);
   U13675 : OAI22_X1 port map( A1 => n16629, A2 => n23562, B1 => n20376, B2 => 
                           n22845, ZN => n3722);
   U13676 : OAI22_X1 port map( A1 => n16623, A2 => n23564, B1 => n20370, B2 => 
                           n22846, ZN => n3728);
   U13677 : OAI22_X1 port map( A1 => n16622, A2 => n23563, B1 => n20369, B2 => 
                           n22846, ZN => n3729);
   U13678 : OAI22_X1 port map( A1 => n16621, A2 => n23562, B1 => n20368, B2 => 
                           n22846, ZN => n3730);
   U13679 : OAI22_X1 port map( A1 => n16620, A2 => n23564, B1 => n20367, B2 => 
                           n22846, ZN => n3731);
   U13680 : OAI22_X1 port map( A1 => n16619, A2 => n23563, B1 => n20366, B2 => 
                           n22846, ZN => n3732);
   U13681 : OAI22_X1 port map( A1 => n16618, A2 => n23562, B1 => n20365, B2 => 
                           n22846, ZN => n3733);
   U13682 : OAI22_X1 port map( A1 => n16617, A2 => n23564, B1 => n20364, B2 => 
                           n22846, ZN => n3734);
   U13683 : OAI22_X1 port map( A1 => n16611, A2 => n23562, B1 => n20358, B2 => 
                           n22847, ZN => n3740);
   U13684 : OAI22_X1 port map( A1 => n16610, A2 => n23562, B1 => n20357, B2 => 
                           n22847, ZN => n3741);
   U13685 : OAI22_X1 port map( A1 => n16609, A2 => n23564, B1 => n20356, B2 => 
                           n22847, ZN => n3742);
   U13686 : OAI22_X1 port map( A1 => n16608, A2 => n23563, B1 => n20355, B2 => 
                           n22847, ZN => n3743);
   U13687 : OAI22_X1 port map( A1 => n16607, A2 => n23562, B1 => n20354, B2 => 
                           n22847, ZN => n3744);
   U13688 : OAI22_X1 port map( A1 => n16606, A2 => n23562, B1 => n20353, B2 => 
                           n22847, ZN => n3745);
   U13689 : OAI22_X1 port map( A1 => n16605, A2 => n23564, B1 => n20352, B2 => 
                           n22847, ZN => n3746);
   U13690 : OAI22_X1 port map( A1 => n16635, A2 => n23582, B1 => n20254, B2 => 
                           n22857, ZN => n3844);
   U13691 : OAI22_X1 port map( A1 => n16634, A2 => n23582, B1 => n20253, B2 => 
                           n22857, ZN => n3845);
   U13692 : OAI22_X1 port map( A1 => n16633, A2 => n23582, B1 => n20252, B2 => 
                           n22857, ZN => n3846);
   U13693 : OAI22_X1 port map( A1 => n16632, A2 => n23582, B1 => n20251, B2 => 
                           n22857, ZN => n3847);
   U13694 : OAI22_X1 port map( A1 => n16631, A2 => n23582, B1 => n20250, B2 => 
                           n22857, ZN => n3848);
   U13695 : OAI22_X1 port map( A1 => n16630, A2 => n23582, B1 => n20249, B2 => 
                           n22857, ZN => n3849);
   U13696 : OAI22_X1 port map( A1 => n16629, A2 => n23582, B1 => n20248, B2 => 
                           n22857, ZN => n3850);
   U13697 : OAI22_X1 port map( A1 => n16623, A2 => n23584, B1 => n20242, B2 => 
                           n22858, ZN => n3856);
   U13698 : OAI22_X1 port map( A1 => n16622, A2 => n23583, B1 => n20241, B2 => 
                           n22858, ZN => n3857);
   U13699 : OAI22_X1 port map( A1 => n16621, A2 => n23582, B1 => n20240, B2 => 
                           n22858, ZN => n3858);
   U13700 : OAI22_X1 port map( A1 => n16620, A2 => n23584, B1 => n20239, B2 => 
                           n22858, ZN => n3859);
   U13701 : OAI22_X1 port map( A1 => n16619, A2 => n23583, B1 => n20238, B2 => 
                           n22858, ZN => n3860);
   U13702 : OAI22_X1 port map( A1 => n16618, A2 => n23582, B1 => n20237, B2 => 
                           n22858, ZN => n3861);
   U13703 : OAI22_X1 port map( A1 => n16617, A2 => n23584, B1 => n20236, B2 => 
                           n22858, ZN => n3862);
   U13704 : OAI22_X1 port map( A1 => n16611, A2 => n23582, B1 => n20230, B2 => 
                           n22859, ZN => n3868);
   U13705 : OAI22_X1 port map( A1 => n16610, A2 => n23582, B1 => n20229, B2 => 
                           n22859, ZN => n3869);
   U13706 : OAI22_X1 port map( A1 => n16609, A2 => n23584, B1 => n20228, B2 => 
                           n22859, ZN => n3870);
   U13707 : OAI22_X1 port map( A1 => n16608, A2 => n23583, B1 => n20227, B2 => 
                           n22859, ZN => n3871);
   U13708 : OAI22_X1 port map( A1 => n16607, A2 => n23582, B1 => n20226, B2 => 
                           n22859, ZN => n3872);
   U13709 : OAI22_X1 port map( A1 => n16606, A2 => n23582, B1 => n20225, B2 => 
                           n22859, ZN => n3873);
   U13710 : OAI22_X1 port map( A1 => n16605, A2 => n23584, B1 => n20224, B2 => 
                           n22859, ZN => n3874);
   U13711 : OAI22_X1 port map( A1 => n16635, A2 => n23532, B1 => n20574, B2 => 
                           n22827, ZN => n3524);
   U13712 : OAI22_X1 port map( A1 => n16634, A2 => n23532, B1 => n20573, B2 => 
                           n22827, ZN => n3525);
   U13713 : OAI22_X1 port map( A1 => n16633, A2 => n23532, B1 => n20572, B2 => 
                           n22827, ZN => n3526);
   U13714 : OAI22_X1 port map( A1 => n16632, A2 => n23532, B1 => n20571, B2 => 
                           n22827, ZN => n3527);
   U13715 : OAI22_X1 port map( A1 => n16631, A2 => n23532, B1 => n20570, B2 => 
                           n22827, ZN => n3528);
   U13716 : OAI22_X1 port map( A1 => n16630, A2 => n23532, B1 => n20569, B2 => 
                           n22827, ZN => n3529);
   U13717 : OAI22_X1 port map( A1 => n16629, A2 => n23532, B1 => n20568, B2 => 
                           n22827, ZN => n3530);
   U13718 : OAI22_X1 port map( A1 => n16623, A2 => n23534, B1 => n20562, B2 => 
                           n22828, ZN => n3536);
   U13719 : OAI22_X1 port map( A1 => n16622, A2 => n23533, B1 => n20561, B2 => 
                           n22828, ZN => n3537);
   U13720 : OAI22_X1 port map( A1 => n16621, A2 => n23532, B1 => n20560, B2 => 
                           n22828, ZN => n3538);
   U13721 : OAI22_X1 port map( A1 => n16620, A2 => n23534, B1 => n20559, B2 => 
                           n22828, ZN => n3539);
   U13722 : OAI22_X1 port map( A1 => n16619, A2 => n23533, B1 => n20558, B2 => 
                           n22828, ZN => n3540);
   U13723 : OAI22_X1 port map( A1 => n16618, A2 => n23532, B1 => n20557, B2 => 
                           n22828, ZN => n3541);
   U13724 : OAI22_X1 port map( A1 => n16617, A2 => n23534, B1 => n20556, B2 => 
                           n22828, ZN => n3542);
   U13725 : OAI22_X1 port map( A1 => n16611, A2 => n23532, B1 => n20550, B2 => 
                           n22829, ZN => n3548);
   U13726 : OAI22_X1 port map( A1 => n16610, A2 => n23532, B1 => n20549, B2 => 
                           n22829, ZN => n3549);
   U13727 : OAI22_X1 port map( A1 => n16609, A2 => n23534, B1 => n20548, B2 => 
                           n22829, ZN => n3550);
   U13728 : OAI22_X1 port map( A1 => n16608, A2 => n23533, B1 => n20547, B2 => 
                           n22829, ZN => n3551);
   U13729 : OAI22_X1 port map( A1 => n16607, A2 => n23532, B1 => n20546, B2 => 
                           n22829, ZN => n3552);
   U13730 : OAI22_X1 port map( A1 => n16606, A2 => n23532, B1 => n20545, B2 => 
                           n22829, ZN => n3553);
   U13731 : OAI22_X1 port map( A1 => n16605, A2 => n23534, B1 => n20544, B2 => 
                           n22829, ZN => n3554);
   U13732 : OAI22_X1 port map( A1 => n16635, A2 => n23552, B1 => n20446, B2 => 
                           n22839, ZN => n3652);
   U13733 : OAI22_X1 port map( A1 => n16634, A2 => n23552, B1 => n20445, B2 => 
                           n22839, ZN => n3653);
   U13734 : OAI22_X1 port map( A1 => n16633, A2 => n23552, B1 => n20444, B2 => 
                           n22839, ZN => n3654);
   U13735 : OAI22_X1 port map( A1 => n16632, A2 => n23552, B1 => n20443, B2 => 
                           n22839, ZN => n3655);
   U13736 : OAI22_X1 port map( A1 => n16631, A2 => n23552, B1 => n20442, B2 => 
                           n22839, ZN => n3656);
   U13737 : OAI22_X1 port map( A1 => n16630, A2 => n23552, B1 => n20441, B2 => 
                           n22839, ZN => n3657);
   U13738 : OAI22_X1 port map( A1 => n16629, A2 => n23552, B1 => n20440, B2 => 
                           n22839, ZN => n3658);
   U13739 : OAI22_X1 port map( A1 => n16623, A2 => n23554, B1 => n20434, B2 => 
                           n22840, ZN => n3664);
   U13740 : OAI22_X1 port map( A1 => n16622, A2 => n23553, B1 => n20433, B2 => 
                           n22840, ZN => n3665);
   U13741 : OAI22_X1 port map( A1 => n16621, A2 => n23552, B1 => n20432, B2 => 
                           n22840, ZN => n3666);
   U13742 : OAI22_X1 port map( A1 => n16620, A2 => n23554, B1 => n20431, B2 => 
                           n22840, ZN => n3667);
   U13743 : OAI22_X1 port map( A1 => n16619, A2 => n23553, B1 => n20430, B2 => 
                           n22840, ZN => n3668);
   U13744 : OAI22_X1 port map( A1 => n16618, A2 => n23552, B1 => n20429, B2 => 
                           n22840, ZN => n3669);
   U13745 : OAI22_X1 port map( A1 => n16617, A2 => n23554, B1 => n20428, B2 => 
                           n22840, ZN => n3670);
   U13746 : OAI22_X1 port map( A1 => n16611, A2 => n23552, B1 => n20422, B2 => 
                           n22841, ZN => n3676);
   U13747 : OAI22_X1 port map( A1 => n16610, A2 => n23552, B1 => n20421, B2 => 
                           n22841, ZN => n3677);
   U13748 : OAI22_X1 port map( A1 => n16609, A2 => n23554, B1 => n20420, B2 => 
                           n22841, ZN => n3678);
   U13749 : OAI22_X1 port map( A1 => n16608, A2 => n23553, B1 => n20419, B2 => 
                           n22841, ZN => n3679);
   U13750 : OAI22_X1 port map( A1 => n16607, A2 => n23552, B1 => n20418, B2 => 
                           n22841, ZN => n3680);
   U13751 : OAI22_X1 port map( A1 => n16606, A2 => n23552, B1 => n20417, B2 => 
                           n22841, ZN => n3681);
   U13752 : OAI22_X1 port map( A1 => n16605, A2 => n23554, B1 => n20416, B2 => 
                           n22841, ZN => n3682);
   U13753 : OAI22_X1 port map( A1 => n16635, A2 => n23572, B1 => n20318, B2 => 
                           n22851, ZN => n3780);
   U13754 : OAI22_X1 port map( A1 => n16634, A2 => n23572, B1 => n20317, B2 => 
                           n22851, ZN => n3781);
   U13755 : OAI22_X1 port map( A1 => n16633, A2 => n23572, B1 => n20316, B2 => 
                           n22851, ZN => n3782);
   U13756 : OAI22_X1 port map( A1 => n16632, A2 => n23572, B1 => n20315, B2 => 
                           n22851, ZN => n3783);
   U13757 : OAI22_X1 port map( A1 => n16631, A2 => n23572, B1 => n20314, B2 => 
                           n22851, ZN => n3784);
   U13758 : OAI22_X1 port map( A1 => n16630, A2 => n23572, B1 => n20313, B2 => 
                           n22851, ZN => n3785);
   U13759 : OAI22_X1 port map( A1 => n16629, A2 => n23572, B1 => n20312, B2 => 
                           n22851, ZN => n3786);
   U13760 : OAI22_X1 port map( A1 => n16623, A2 => n23574, B1 => n20306, B2 => 
                           n22852, ZN => n3792);
   U13761 : OAI22_X1 port map( A1 => n16622, A2 => n23573, B1 => n20305, B2 => 
                           n22852, ZN => n3793);
   U13762 : OAI22_X1 port map( A1 => n16621, A2 => n23572, B1 => n20304, B2 => 
                           n22852, ZN => n3794);
   U13763 : OAI22_X1 port map( A1 => n16620, A2 => n23574, B1 => n20303, B2 => 
                           n22852, ZN => n3795);
   U13764 : OAI22_X1 port map( A1 => n16619, A2 => n23573, B1 => n20302, B2 => 
                           n22852, ZN => n3796);
   U13765 : OAI22_X1 port map( A1 => n16618, A2 => n23572, B1 => n20301, B2 => 
                           n22852, ZN => n3797);
   U13766 : OAI22_X1 port map( A1 => n16617, A2 => n23574, B1 => n20300, B2 => 
                           n22852, ZN => n3798);
   U13767 : OAI22_X1 port map( A1 => n16611, A2 => n23572, B1 => n20294, B2 => 
                           n22853, ZN => n3804);
   U13768 : OAI22_X1 port map( A1 => n16610, A2 => n23572, B1 => n20293, B2 => 
                           n22853, ZN => n3805);
   U13769 : OAI22_X1 port map( A1 => n16609, A2 => n23574, B1 => n20292, B2 => 
                           n22853, ZN => n3806);
   U13770 : OAI22_X1 port map( A1 => n16608, A2 => n23573, B1 => n20291, B2 => 
                           n22853, ZN => n3807);
   U13771 : OAI22_X1 port map( A1 => n16607, A2 => n23572, B1 => n20290, B2 => 
                           n22853, ZN => n3808);
   U13772 : OAI22_X1 port map( A1 => n16606, A2 => n23572, B1 => n20289, B2 => 
                           n22853, ZN => n3809);
   U13773 : OAI22_X1 port map( A1 => n16605, A2 => n23574, B1 => n20288, B2 => 
                           n22853, ZN => n3810);
   U13774 : OAI22_X1 port map( A1 => n16636, A2 => n23582, B1 => n20255, B2 => 
                           n22857, ZN => n3843);
   U13775 : OAI22_X1 port map( A1 => n16628, A2 => n23582, B1 => n20247, B2 => 
                           n22860, ZN => n3851);
   U13776 : OAI22_X1 port map( A1 => n16627, A2 => n23582, B1 => n20246, B2 => 
                           n22858, ZN => n3852);
   U13777 : OAI22_X1 port map( A1 => n16626, A2 => n23582, B1 => n20245, B2 => 
                           n22858, ZN => n3853);
   U13778 : OAI22_X1 port map( A1 => n16625, A2 => n23582, B1 => n20244, B2 => 
                           n22858, ZN => n3854);
   U13779 : OAI22_X1 port map( A1 => n16624, A2 => n23583, B1 => n20243, B2 => 
                           n22858, ZN => n3855);
   U13780 : OAI22_X1 port map( A1 => n16616, A2 => n23582, B1 => n20235, B2 => 
                           n22858, ZN => n3863);
   U13781 : OAI22_X1 port map( A1 => n16615, A2 => n23584, B1 => n20234, B2 => 
                           n22859, ZN => n3864);
   U13782 : OAI22_X1 port map( A1 => n16614, A2 => n23583, B1 => n20233, B2 => 
                           n22859, ZN => n3865);
   U13783 : OAI22_X1 port map( A1 => n16613, A2 => n23582, B1 => n20232, B2 => 
                           n22859, ZN => n3866);
   U13784 : OAI22_X1 port map( A1 => n16612, A2 => n23583, B1 => n20231, B2 => 
                           n22859, ZN => n3867);
   U13785 : OAI22_X1 port map( A1 => n16604, A2 => n23582, B1 => n20223, B2 => 
                           n22859, ZN => n3875);
   U13786 : OAI22_X1 port map( A1 => n16603, A2 => n23584, B1 => n20222, B2 => 
                           n22860, ZN => n3876);
   U13787 : OAI22_X1 port map( A1 => n16602, A2 => n23584, B1 => n20221, B2 => 
                           n22860, ZN => n3877);
   U13788 : OAI22_X1 port map( A1 => n16601, A2 => n23583, B1 => n20220, B2 => 
                           n22860, ZN => n3878);
   U13789 : OAI22_X1 port map( A1 => n16636, A2 => n23532, B1 => n20575, B2 => 
                           n22827, ZN => n3523);
   U13790 : OAI22_X1 port map( A1 => n16628, A2 => n23532, B1 => n20567, B2 => 
                           n22830, ZN => n3531);
   U13791 : OAI22_X1 port map( A1 => n16627, A2 => n23532, B1 => n20566, B2 => 
                           n22828, ZN => n3532);
   U13792 : OAI22_X1 port map( A1 => n16626, A2 => n23532, B1 => n20565, B2 => 
                           n22828, ZN => n3533);
   U13793 : OAI22_X1 port map( A1 => n16625, A2 => n23532, B1 => n20564, B2 => 
                           n22828, ZN => n3534);
   U13794 : OAI22_X1 port map( A1 => n16624, A2 => n23533, B1 => n20563, B2 => 
                           n22828, ZN => n3535);
   U13795 : OAI22_X1 port map( A1 => n16616, A2 => n23532, B1 => n20555, B2 => 
                           n22828, ZN => n3543);
   U13796 : OAI22_X1 port map( A1 => n16615, A2 => n23534, B1 => n20554, B2 => 
                           n22829, ZN => n3544);
   U13797 : OAI22_X1 port map( A1 => n16614, A2 => n23533, B1 => n20553, B2 => 
                           n22829, ZN => n3545);
   U13798 : OAI22_X1 port map( A1 => n16613, A2 => n23532, B1 => n20552, B2 => 
                           n22829, ZN => n3546);
   U13799 : OAI22_X1 port map( A1 => n16612, A2 => n23533, B1 => n20551, B2 => 
                           n22829, ZN => n3547);
   U13800 : OAI22_X1 port map( A1 => n16604, A2 => n23532, B1 => n20543, B2 => 
                           n22829, ZN => n3555);
   U13801 : OAI22_X1 port map( A1 => n16603, A2 => n23534, B1 => n20542, B2 => 
                           n22830, ZN => n3556);
   U13802 : OAI22_X1 port map( A1 => n16602, A2 => n23534, B1 => n20541, B2 => 
                           n22830, ZN => n3557);
   U13803 : OAI22_X1 port map( A1 => n16601, A2 => n23533, B1 => n20540, B2 => 
                           n22830, ZN => n3558);
   U13804 : OAI22_X1 port map( A1 => n16636, A2 => n23552, B1 => n20447, B2 => 
                           n22839, ZN => n3651);
   U13805 : OAI22_X1 port map( A1 => n16628, A2 => n23552, B1 => n20439, B2 => 
                           n22842, ZN => n3659);
   U13806 : OAI22_X1 port map( A1 => n16627, A2 => n23552, B1 => n20438, B2 => 
                           n22840, ZN => n3660);
   U13807 : OAI22_X1 port map( A1 => n16626, A2 => n23552, B1 => n20437, B2 => 
                           n22840, ZN => n3661);
   U13808 : OAI22_X1 port map( A1 => n16625, A2 => n23552, B1 => n20436, B2 => 
                           n22840, ZN => n3662);
   U13809 : OAI22_X1 port map( A1 => n16624, A2 => n23553, B1 => n20435, B2 => 
                           n22840, ZN => n3663);
   U13810 : OAI22_X1 port map( A1 => n16616, A2 => n23552, B1 => n20427, B2 => 
                           n22840, ZN => n3671);
   U13811 : OAI22_X1 port map( A1 => n16615, A2 => n23554, B1 => n20426, B2 => 
                           n22841, ZN => n3672);
   U13812 : OAI22_X1 port map( A1 => n16614, A2 => n23553, B1 => n20425, B2 => 
                           n22841, ZN => n3673);
   U13813 : OAI22_X1 port map( A1 => n16613, A2 => n23552, B1 => n20424, B2 => 
                           n22841, ZN => n3674);
   U13814 : OAI22_X1 port map( A1 => n16612, A2 => n23553, B1 => n20423, B2 => 
                           n22841, ZN => n3675);
   U13815 : OAI22_X1 port map( A1 => n16604, A2 => n23552, B1 => n20415, B2 => 
                           n22841, ZN => n3683);
   U13816 : OAI22_X1 port map( A1 => n16603, A2 => n23554, B1 => n20414, B2 => 
                           n22842, ZN => n3684);
   U13817 : OAI22_X1 port map( A1 => n16602, A2 => n23554, B1 => n20413, B2 => 
                           n22842, ZN => n3685);
   U13818 : OAI22_X1 port map( A1 => n16601, A2 => n23553, B1 => n20412, B2 => 
                           n22842, ZN => n3686);
   U13819 : OAI22_X1 port map( A1 => n16636, A2 => n23542, B1 => n20511, B2 => 
                           n22833, ZN => n3587);
   U13820 : OAI22_X1 port map( A1 => n16628, A2 => n23542, B1 => n20503, B2 => 
                           n22836, ZN => n3595);
   U13821 : OAI22_X1 port map( A1 => n16627, A2 => n23542, B1 => n20502, B2 => 
                           n22834, ZN => n3596);
   U13822 : OAI22_X1 port map( A1 => n16626, A2 => n23542, B1 => n20501, B2 => 
                           n22834, ZN => n3597);
   U13823 : OAI22_X1 port map( A1 => n16625, A2 => n23542, B1 => n20500, B2 => 
                           n22834, ZN => n3598);
   U13824 : OAI22_X1 port map( A1 => n16624, A2 => n23543, B1 => n20499, B2 => 
                           n22834, ZN => n3599);
   U13825 : OAI22_X1 port map( A1 => n16616, A2 => n23542, B1 => n20491, B2 => 
                           n22834, ZN => n3607);
   U13826 : OAI22_X1 port map( A1 => n16615, A2 => n23544, B1 => n20490, B2 => 
                           n22835, ZN => n3608);
   U13827 : OAI22_X1 port map( A1 => n16614, A2 => n23543, B1 => n20489, B2 => 
                           n22835, ZN => n3609);
   U13828 : OAI22_X1 port map( A1 => n16613, A2 => n23542, B1 => n20488, B2 => 
                           n22835, ZN => n3610);
   U13829 : OAI22_X1 port map( A1 => n16612, A2 => n23543, B1 => n20487, B2 => 
                           n22835, ZN => n3611);
   U13830 : OAI22_X1 port map( A1 => n16604, A2 => n23542, B1 => n20479, B2 => 
                           n22835, ZN => n3619);
   U13831 : OAI22_X1 port map( A1 => n16603, A2 => n23544, B1 => n20478, B2 => 
                           n22836, ZN => n3620);
   U13832 : OAI22_X1 port map( A1 => n16602, A2 => n23544, B1 => n20477, B2 => 
                           n22836, ZN => n3621);
   U13833 : OAI22_X1 port map( A1 => n16601, A2 => n23543, B1 => n20476, B2 => 
                           n22836, ZN => n3622);
   U13834 : OAI22_X1 port map( A1 => n16636, A2 => n23522, B1 => n20639, B2 => 
                           n22821, ZN => n3459);
   U13835 : OAI22_X1 port map( A1 => n16628, A2 => n23522, B1 => n20631, B2 => 
                           n22824, ZN => n3467);
   U13836 : OAI22_X1 port map( A1 => n16627, A2 => n23522, B1 => n20630, B2 => 
                           n22822, ZN => n3468);
   U13837 : OAI22_X1 port map( A1 => n16626, A2 => n23522, B1 => n20629, B2 => 
                           n22822, ZN => n3469);
   U13838 : OAI22_X1 port map( A1 => n16625, A2 => n23522, B1 => n20628, B2 => 
                           n22822, ZN => n3470);
   U13839 : OAI22_X1 port map( A1 => n16624, A2 => n23523, B1 => n20627, B2 => 
                           n22822, ZN => n3471);
   U13840 : OAI22_X1 port map( A1 => n16616, A2 => n23522, B1 => n20619, B2 => 
                           n22822, ZN => n3479);
   U13841 : OAI22_X1 port map( A1 => n16615, A2 => n23524, B1 => n20618, B2 => 
                           n22823, ZN => n3480);
   U13842 : OAI22_X1 port map( A1 => n16614, A2 => n23523, B1 => n20617, B2 => 
                           n22823, ZN => n3481);
   U13843 : OAI22_X1 port map( A1 => n16613, A2 => n23522, B1 => n20616, B2 => 
                           n22823, ZN => n3482);
   U13844 : OAI22_X1 port map( A1 => n16612, A2 => n23523, B1 => n20615, B2 => 
                           n22823, ZN => n3483);
   U13845 : OAI22_X1 port map( A1 => n16604, A2 => n23522, B1 => n20607, B2 => 
                           n22823, ZN => n3491);
   U13846 : OAI22_X1 port map( A1 => n16603, A2 => n23524, B1 => n20606, B2 => 
                           n22824, ZN => n3492);
   U13847 : OAI22_X1 port map( A1 => n16602, A2 => n23524, B1 => n20605, B2 => 
                           n22824, ZN => n3493);
   U13848 : OAI22_X1 port map( A1 => n16601, A2 => n23523, B1 => n20604, B2 => 
                           n22824, ZN => n3494);
   U13849 : OAI22_X1 port map( A1 => n16636, A2 => n23562, B1 => n20383, B2 => 
                           n22845, ZN => n3715);
   U13850 : OAI22_X1 port map( A1 => n16628, A2 => n23562, B1 => n20375, B2 => 
                           n22848, ZN => n3723);
   U13851 : OAI22_X1 port map( A1 => n16627, A2 => n23562, B1 => n20374, B2 => 
                           n22846, ZN => n3724);
   U13852 : OAI22_X1 port map( A1 => n16626, A2 => n23562, B1 => n20373, B2 => 
                           n22846, ZN => n3725);
   U13853 : OAI22_X1 port map( A1 => n16625, A2 => n23562, B1 => n20372, B2 => 
                           n22846, ZN => n3726);
   U13854 : OAI22_X1 port map( A1 => n16624, A2 => n23563, B1 => n20371, B2 => 
                           n22846, ZN => n3727);
   U13855 : OAI22_X1 port map( A1 => n16616, A2 => n23562, B1 => n20363, B2 => 
                           n22846, ZN => n3735);
   U13856 : OAI22_X1 port map( A1 => n16615, A2 => n23564, B1 => n20362, B2 => 
                           n22847, ZN => n3736);
   U13857 : OAI22_X1 port map( A1 => n16614, A2 => n23563, B1 => n20361, B2 => 
                           n22847, ZN => n3737);
   U13858 : OAI22_X1 port map( A1 => n16613, A2 => n23562, B1 => n20360, B2 => 
                           n22847, ZN => n3738);
   U13859 : OAI22_X1 port map( A1 => n16612, A2 => n23563, B1 => n20359, B2 => 
                           n22847, ZN => n3739);
   U13860 : OAI22_X1 port map( A1 => n16604, A2 => n23562, B1 => n20351, B2 => 
                           n22847, ZN => n3747);
   U13861 : OAI22_X1 port map( A1 => n16603, A2 => n23564, B1 => n20350, B2 => 
                           n22848, ZN => n3748);
   U13862 : OAI22_X1 port map( A1 => n16602, A2 => n23564, B1 => n20349, B2 => 
                           n22848, ZN => n3749);
   U13863 : OAI22_X1 port map( A1 => n16601, A2 => n23563, B1 => n20348, B2 => 
                           n22848, ZN => n3750);
   U13864 : OAI22_X1 port map( A1 => n16636, A2 => n23572, B1 => n20319, B2 => 
                           n22851, ZN => n3779);
   U13865 : OAI22_X1 port map( A1 => n16628, A2 => n23572, B1 => n20311, B2 => 
                           n22854, ZN => n3787);
   U13866 : OAI22_X1 port map( A1 => n16627, A2 => n23572, B1 => n20310, B2 => 
                           n22852, ZN => n3788);
   U13867 : OAI22_X1 port map( A1 => n16626, A2 => n23572, B1 => n20309, B2 => 
                           n22852, ZN => n3789);
   U13868 : OAI22_X1 port map( A1 => n16625, A2 => n23572, B1 => n20308, B2 => 
                           n22852, ZN => n3790);
   U13869 : OAI22_X1 port map( A1 => n16624, A2 => n23573, B1 => n20307, B2 => 
                           n22852, ZN => n3791);
   U13870 : OAI22_X1 port map( A1 => n16616, A2 => n23572, B1 => n20299, B2 => 
                           n22852, ZN => n3799);
   U13871 : OAI22_X1 port map( A1 => n16615, A2 => n23574, B1 => n20298, B2 => 
                           n22853, ZN => n3800);
   U13872 : OAI22_X1 port map( A1 => n16614, A2 => n23573, B1 => n20297, B2 => 
                           n22853, ZN => n3801);
   U13873 : OAI22_X1 port map( A1 => n16613, A2 => n23572, B1 => n20296, B2 => 
                           n22853, ZN => n3802);
   U13874 : OAI22_X1 port map( A1 => n16612, A2 => n23573, B1 => n20295, B2 => 
                           n22853, ZN => n3803);
   U13875 : OAI22_X1 port map( A1 => n16604, A2 => n23572, B1 => n20287, B2 => 
                           n22853, ZN => n3811);
   U13876 : OAI22_X1 port map( A1 => n16603, A2 => n23574, B1 => n20286, B2 => 
                           n22854, ZN => n3812);
   U13877 : OAI22_X1 port map( A1 => n16602, A2 => n23574, B1 => n20285, B2 => 
                           n22854, ZN => n3813);
   U13878 : OAI22_X1 port map( A1 => n16601, A2 => n23573, B1 => n20284, B2 => 
                           n22854, ZN => n3814);
   U13879 : AOI221_X1 port map( B1 => n23833, B2 => n21766, C1 => n23826, C2 =>
                           n22291, A => n16542, ZN => n16538);
   U13880 : OAI22_X1 port map( A1 => n18780, A2 => n23286, B1 => n18908, B2 => 
                           n23298, ZN => n16542);
   U13881 : AOI221_X1 port map( B1 => n23865, B2 => n21285, C1 => n23849, C2 =>
                           n21842, A => n16541, ZN => n16539);
   U13882 : OAI22_X1 port map( A1 => n18972, A2 => n23309, B1 => n19100, B2 => 
                           n23321, ZN => n16541);
   U13883 : AOI221_X1 port map( B1 => n23865, B2 => n21265, C1 => n23849, C2 =>
                           n21750, A => n16518, ZN => n16517);
   U13884 : OAI22_X1 port map( A1 => n18940, A2 => n23309, B1 => n19068, B2 => 
                           n23321, ZN => n16518);
   U13885 : AOI221_X1 port map( B1 => n23865, B2 => n21242, C1 => n23849, C2 =>
                           n21727, A => n16497, ZN => n16496);
   U13886 : OAI22_X1 port map( A1 => n19003, A2 => n23309, B1 => n19131, B2 => 
                           n23321, ZN => n16497);
   U13887 : AOI221_X1 port map( B1 => n23865, B2 => n21264, C1 => n23849, C2 =>
                           n21749, A => n16476, ZN => n16475);
   U13888 : OAI22_X1 port map( A1 => n18941, A2 => n23309, B1 => n19069, B2 => 
                           n23321, ZN => n16476);
   U13889 : AOI221_X1 port map( B1 => n23865, B2 => n21263, C1 => n23849, C2 =>
                           n21748, A => n16455, ZN => n16454);
   U13890 : OAI22_X1 port map( A1 => n19002, A2 => n23309, B1 => n19130, B2 => 
                           n23321, ZN => n16455);
   U13891 : AOI221_X1 port map( B1 => n23866, B2 => n21224, C1 => n23850, C2 =>
                           n21709, A => n16434, ZN => n16433);
   U13892 : OAI22_X1 port map( A1 => n18942, A2 => n23309, B1 => n19070, B2 => 
                           n23321, ZN => n16434);
   U13893 : AOI221_X1 port map( B1 => n23866, B2 => n21262, C1 => n23850, C2 =>
                           n21747, A => n16413, ZN => n16412);
   U13894 : OAI22_X1 port map( A1 => n19001, A2 => n23310, B1 => n19129, B2 => 
                           n23322, ZN => n16413);
   U13895 : AOI221_X1 port map( B1 => n23866, B2 => n21261, C1 => n23850, C2 =>
                           n21746, A => n16392, ZN => n16391);
   U13896 : OAI22_X1 port map( A1 => n18943, A2 => n23310, B1 => n19071, B2 => 
                           n23322, ZN => n16392);
   U13897 : AOI221_X1 port map( B1 => n23866, B2 => n21223, C1 => n23850, C2 =>
                           n21708, A => n16371, ZN => n16370);
   U13898 : OAI22_X1 port map( A1 => n19000, A2 => n23310, B1 => n19128, B2 => 
                           n23322, ZN => n16371);
   U13899 : AOI221_X1 port map( B1 => n23866, B2 => n21243, C1 => n23850, C2 =>
                           n21745, A => n16350, ZN => n16349);
   U13900 : OAI22_X1 port map( A1 => n18944, A2 => n23310, B1 => n19072, B2 => 
                           n23322, ZN => n16350);
   U13901 : AOI221_X1 port map( B1 => n23866, B2 => n21260, C1 => n23850, C2 =>
                           n21744, A => n16329, ZN => n16328);
   U13902 : OAI22_X1 port map( A1 => n18999, A2 => n23310, B1 => n19127, B2 => 
                           n23322, ZN => n16329);
   U13903 : AOI221_X1 port map( B1 => n23866, B2 => n21222, C1 => n23850, C2 =>
                           n21707, A => n16308, ZN => n16307);
   U13904 : OAI22_X1 port map( A1 => n18945, A2 => n23310, B1 => n19073, B2 => 
                           n23322, ZN => n16308);
   U13905 : AOI221_X1 port map( B1 => n23833, B2 => n21825, C1 => n23826, C2 =>
                           n22057, A => n16519, ZN => n16516);
   U13906 : OAI22_X1 port map( A1 => n18748, A2 => n23286, B1 => n18876, B2 => 
                           n23298, ZN => n16519);
   U13907 : AOI221_X1 port map( B1 => n23833, B2 => n21824, C1 => n23826, C2 =>
                           n22183, A => n16498, ZN => n16495);
   U13908 : OAI22_X1 port map( A1 => n18811, A2 => n23286, B1 => n18939, B2 => 
                           n23298, ZN => n16498);
   U13909 : AOI221_X1 port map( B1 => n23833, B2 => n21823, C1 => n23826, C2 =>
                           n22182, A => n16477, ZN => n16474);
   U13910 : OAI22_X1 port map( A1 => n18749, A2 => n23286, B1 => n18877, B2 => 
                           n23298, ZN => n16477);
   U13911 : AOI221_X1 port map( B1 => n23833, B2 => n21822, C1 => n23825, C2 =>
                           n22181, A => n16456, ZN => n16453);
   U13912 : OAI22_X1 port map( A1 => n18810, A2 => n23286, B1 => n18938, B2 => 
                           n23298, ZN => n16456);
   U13913 : AOI221_X1 port map( B1 => n23834, B2 => n21821, C1 => n23825, C2 =>
                           n22056, A => n16435, ZN => n16432);
   U13914 : OAI22_X1 port map( A1 => n18750, A2 => n23286, B1 => n18878, B2 => 
                           n23298, ZN => n16435);
   U13915 : AOI221_X1 port map( B1 => n23834, B2 => n21820, C1 => n23825, C2 =>
                           n22180, A => n16414, ZN => n16411);
   U13916 : OAI22_X1 port map( A1 => n18809, A2 => n23287, B1 => n18937, B2 => 
                           n23299, ZN => n16414);
   U13917 : AOI221_X1 port map( B1 => n23834, B2 => n21819, C1 => n23825, C2 =>
                           n22179, A => n16393, ZN => n16390);
   U13918 : OAI22_X1 port map( A1 => n18751, A2 => n23287, B1 => n18879, B2 => 
                           n23299, ZN => n16393);
   U13919 : AOI221_X1 port map( B1 => n23834, B2 => n21818, C1 => n23825, C2 =>
                           n22178, A => n16372, ZN => n16369);
   U13920 : OAI22_X1 port map( A1 => n18808, A2 => n23287, B1 => n18936, B2 => 
                           n23299, ZN => n16372);
   U13921 : AOI221_X1 port map( B1 => n23834, B2 => n21817, C1 => n23825, C2 =>
                           n22036, A => n16351, ZN => n16348);
   U13922 : OAI22_X1 port map( A1 => n18752, A2 => n23287, B1 => n18880, B2 => 
                           n23299, ZN => n16351);
   U13923 : AOI221_X1 port map( B1 => n23834, B2 => n21816, C1 => n23824, C2 =>
                           n22177, A => n16330, ZN => n16327);
   U13924 : OAI22_X1 port map( A1 => n18807, A2 => n23287, B1 => n18935, B2 => 
                           n23299, ZN => n16330);
   U13925 : AOI221_X1 port map( B1 => n23834, B2 => n21815, C1 => n23824, C2 =>
                           n22055, A => n16309, ZN => n16306);
   U13926 : OAI22_X1 port map( A1 => n18753, A2 => n23287, B1 => n18881, B2 => 
                           n23299, ZN => n16309);
   U13927 : AOI221_X1 port map( B1 => n23833, B2 => n22373, C1 => n23826, C2 =>
                           n22336, A => n16523, ZN => n16520);
   U13928 : OAI22_X1 port map( A1 => n19260, A2 => n23286, B1 => n19388, B2 => 
                           n23298, ZN => n16523);
   U13929 : AOI221_X1 port map( B1 => n23833, B2 => n22416, C1 => n23826, C2 =>
                           n22371, A => n16502, ZN => n16499);
   U13930 : OAI22_X1 port map( A1 => n19323, A2 => n23286, B1 => n19451, B2 => 
                           n23298, ZN => n16502);
   U13931 : AOI221_X1 port map( B1 => n23833, B2 => n22374, C1 => n23826, C2 =>
                           n22397, A => n16481, ZN => n16478);
   U13932 : OAI22_X1 port map( A1 => n19261, A2 => n23286, B1 => n19389, B2 => 
                           n23298, ZN => n16481);
   U13933 : AOI221_X1 port map( B1 => n23833, B2 => n22415, C1 => n23825, C2 =>
                           n22410, A => n16460, ZN => n16457);
   U13934 : OAI22_X1 port map( A1 => n19322, A2 => n23286, B1 => n19450, B2 => 
                           n23298, ZN => n16460);
   U13935 : AOI221_X1 port map( B1 => n23833, B2 => n22375, C1 => n23825, C2 =>
                           n22337, A => n16439, ZN => n16436);
   U13936 : OAI22_X1 port map( A1 => n19262, A2 => n23286, B1 => n19390, B2 => 
                           n23298, ZN => n16439);
   U13937 : AOI221_X1 port map( B1 => n23834, B2 => n22414, C1 => n23825, C2 =>
                           n22370, A => n16418, ZN => n16415);
   U13938 : OAI22_X1 port map( A1 => n19321, A2 => n23287, B1 => n19449, B2 => 
                           n23299, ZN => n16418);
   U13939 : AOI221_X1 port map( B1 => n23834, B2 => n22376, C1 => n23825, C2 =>
                           n22358, A => n16397, ZN => n16394);
   U13940 : OAI22_X1 port map( A1 => n19263, A2 => n23287, B1 => n19391, B2 => 
                           n23299, ZN => n16397);
   U13941 : AOI221_X1 port map( B1 => n23834, B2 => n22413, C1 => n23825, C2 =>
                           n22401, A => n16376, ZN => n16373);
   U13942 : OAI22_X1 port map( A1 => n19320, A2 => n23287, B1 => n19448, B2 => 
                           n23299, ZN => n16376);
   U13943 : AOI221_X1 port map( B1 => n23834, B2 => n22367, C1 => n23825, C2 =>
                           n22338, A => n16355, ZN => n16352);
   U13944 : OAI22_X1 port map( A1 => n19264, A2 => n23287, B1 => n19392, B2 => 
                           n23299, ZN => n16355);
   U13945 : AOI221_X1 port map( B1 => n23834, B2 => n22412, C1 => n23824, C2 =>
                           n22369, A => n16334, ZN => n16331);
   U13946 : OAI22_X1 port map( A1 => n19319, A2 => n23287, B1 => n19447, B2 => 
                           n23299, ZN => n16334);
   U13947 : AOI221_X1 port map( B1 => n23834, B2 => n22311, C1 => n23824, C2 =>
                           n22292, A => n16313, ZN => n16310);
   U13948 : OAI22_X1 port map( A1 => n19265, A2 => n23287, B1 => n19393, B2 => 
                           n23299, ZN => n16313);
   U13949 : AOI221_X1 port map( B1 => n23833, B2 => n22372, C1 => n23826, C2 =>
                           n22290, A => n16549, ZN => n16543);
   U13950 : OAI22_X1 port map( A1 => n19292, A2 => n23286, B1 => n19420, B2 => 
                           n23298, ZN => n16549);
   U13951 : AOI221_X1 port map( B1 => n23865, B2 => n21286, C1 => n23849, C2 =>
                           n21840, A => n16546, ZN => n16544);
   U13952 : OAI22_X1 port map( A1 => n19484, A2 => n23309, B1 => n19612, B2 => 
                           n23321, ZN => n16546);
   U13953 : AOI221_X1 port map( B1 => n23865, B2 => n21206, C1 => n23849, C2 =>
                           n21635, A => n16522, ZN => n16521);
   U13954 : OAI22_X1 port map( A1 => n19452, A2 => n23309, B1 => n19580, B2 => 
                           n23321, ZN => n16522);
   U13955 : AOI221_X1 port map( B1 => n23865, B2 => n21203, C1 => n23849, C2 =>
                           n21632, A => n16501, ZN => n16500);
   U13956 : OAI22_X1 port map( A1 => n19515, A2 => n23309, B1 => n19643, B2 => 
                           n23321, ZN => n16501);
   U13957 : AOI221_X1 port map( B1 => n23865, B2 => n21205, C1 => n23849, C2 =>
                           n21634, A => n16480, ZN => n16479);
   U13958 : OAI22_X1 port map( A1 => n19453, A2 => n23309, B1 => n19581, B2 => 
                           n23321, ZN => n16480);
   U13959 : AOI221_X1 port map( B1 => n23865, B2 => n21204, C1 => n23849, C2 =>
                           n21633, A => n16459, ZN => n16458);
   U13960 : OAI22_X1 port map( A1 => n19514, A2 => n23309, B1 => n19642, B2 => 
                           n23321, ZN => n16459);
   U13961 : AOI221_X1 port map( B1 => n23865, B2 => n21181, C1 => n23849, C2 =>
                           n21593, A => n16438, ZN => n16437);
   U13962 : OAI22_X1 port map( A1 => n19454, A2 => n23309, B1 => n19582, B2 => 
                           n23321, ZN => n16438);
   U13963 : AOI221_X1 port map( B1 => n23866, B2 => n21202, C1 => n23850, C2 =>
                           n21630, A => n16417, ZN => n16416);
   U13964 : OAI22_X1 port map( A1 => n19513, A2 => n23310, B1 => n19641, B2 => 
                           n23322, ZN => n16417);
   U13965 : AOI221_X1 port map( B1 => n23866, B2 => n21173, C1 => n23850, C2 =>
                           n21629, A => n16396, ZN => n16395);
   U13966 : OAI22_X1 port map( A1 => n19455, A2 => n23310, B1 => n19583, B2 => 
                           n23322, ZN => n16396);
   U13967 : AOI221_X1 port map( B1 => n23866, B2 => n21180, C1 => n23850, C2 =>
                           n21592, A => n16375, ZN => n16374);
   U13968 : OAI22_X1 port map( A1 => n19512, A2 => n23310, B1 => n19640, B2 => 
                           n23322, ZN => n16375);
   U13969 : AOI221_X1 port map( B1 => n23866, B2 => n21201, C1 => n23850, C2 =>
                           n21628, A => n16354, ZN => n16353);
   U13970 : OAI22_X1 port map( A1 => n19456, A2 => n23310, B1 => n19584, B2 => 
                           n23322, ZN => n16354);
   U13971 : AOI221_X1 port map( B1 => n23866, B2 => n21200, C1 => n23850, C2 =>
                           n21627, A => n16333, ZN => n16332);
   U13972 : OAI22_X1 port map( A1 => n19511, A2 => n23310, B1 => n19639, B2 => 
                           n23322, ZN => n16333);
   U13973 : AOI221_X1 port map( B1 => n23866, B2 => n21179, C1 => n23850, C2 =>
                           n21591, A => n16312, ZN => n16311);
   U13974 : OAI22_X1 port map( A1 => n19457, A2 => n23310, B1 => n19585, B2 => 
                           n23322, ZN => n16312);
   U13975 : OAI22_X1 port map( A1 => n16635, A2 => n23602, B1 => n20126, B2 => 
                           n22869, ZN => n3972);
   U13976 : OAI22_X1 port map( A1 => n16634, A2 => n23602, B1 => n20125, B2 => 
                           n22869, ZN => n3973);
   U13977 : OAI22_X1 port map( A1 => n16633, A2 => n23602, B1 => n20124, B2 => 
                           n22869, ZN => n3974);
   U13978 : OAI22_X1 port map( A1 => n16632, A2 => n23602, B1 => n20123, B2 => 
                           n22869, ZN => n3975);
   U13979 : OAI22_X1 port map( A1 => n16631, A2 => n23602, B1 => n20122, B2 => 
                           n22869, ZN => n3976);
   U13980 : OAI22_X1 port map( A1 => n16630, A2 => n23602, B1 => n20121, B2 => 
                           n22869, ZN => n3977);
   U13981 : OAI22_X1 port map( A1 => n16629, A2 => n23602, B1 => n20120, B2 => 
                           n22869, ZN => n3978);
   U13982 : OAI22_X1 port map( A1 => n16623, A2 => n23604, B1 => n20114, B2 => 
                           n22870, ZN => n3984);
   U13983 : OAI22_X1 port map( A1 => n16622, A2 => n23603, B1 => n20113, B2 => 
                           n22870, ZN => n3985);
   U13984 : OAI22_X1 port map( A1 => n16621, A2 => n23602, B1 => n20112, B2 => 
                           n22870, ZN => n3986);
   U13985 : OAI22_X1 port map( A1 => n16620, A2 => n23604, B1 => n20111, B2 => 
                           n22870, ZN => n3987);
   U13986 : OAI22_X1 port map( A1 => n16619, A2 => n23603, B1 => n20110, B2 => 
                           n22870, ZN => n3988);
   U13987 : OAI22_X1 port map( A1 => n16618, A2 => n23602, B1 => n20109, B2 => 
                           n22870, ZN => n3989);
   U13988 : OAI22_X1 port map( A1 => n16617, A2 => n23604, B1 => n20108, B2 => 
                           n22870, ZN => n3990);
   U13989 : OAI22_X1 port map( A1 => n16611, A2 => n23602, B1 => n20102, B2 => 
                           n22871, ZN => n3996);
   U13990 : OAI22_X1 port map( A1 => n16610, A2 => n23602, B1 => n20101, B2 => 
                           n22871, ZN => n3997);
   U13991 : OAI22_X1 port map( A1 => n16609, A2 => n23604, B1 => n20100, B2 => 
                           n22871, ZN => n3998);
   U13992 : OAI22_X1 port map( A1 => n16608, A2 => n23603, B1 => n20099, B2 => 
                           n22871, ZN => n3999);
   U13993 : OAI22_X1 port map( A1 => n16607, A2 => n23602, B1 => n20098, B2 => 
                           n22871, ZN => n4000);
   U13994 : OAI22_X1 port map( A1 => n16606, A2 => n23602, B1 => n20097, B2 => 
                           n22871, ZN => n4001);
   U13995 : OAI22_X1 port map( A1 => n16605, A2 => n23604, B1 => n20096, B2 => 
                           n22871, ZN => n4002);
   U13996 : OAI22_X1 port map( A1 => n16635, A2 => n23622, B1 => n19998, B2 => 
                           n22881, ZN => n4100);
   U13997 : OAI22_X1 port map( A1 => n16634, A2 => n23622, B1 => n19997, B2 => 
                           n22881, ZN => n4101);
   U13998 : OAI22_X1 port map( A1 => n16633, A2 => n23622, B1 => n19996, B2 => 
                           n22881, ZN => n4102);
   U13999 : OAI22_X1 port map( A1 => n16632, A2 => n23622, B1 => n19995, B2 => 
                           n22881, ZN => n4103);
   U14000 : OAI22_X1 port map( A1 => n16631, A2 => n23622, B1 => n19994, B2 => 
                           n22881, ZN => n4104);
   U14001 : OAI22_X1 port map( A1 => n16630, A2 => n23622, B1 => n19993, B2 => 
                           n22881, ZN => n4105);
   U14002 : OAI22_X1 port map( A1 => n16629, A2 => n23622, B1 => n19992, B2 => 
                           n22881, ZN => n4106);
   U14003 : OAI22_X1 port map( A1 => n16623, A2 => n23624, B1 => n19986, B2 => 
                           n22882, ZN => n4112);
   U14004 : OAI22_X1 port map( A1 => n16622, A2 => n23623, B1 => n19985, B2 => 
                           n22882, ZN => n4113);
   U14005 : OAI22_X1 port map( A1 => n16621, A2 => n23622, B1 => n19984, B2 => 
                           n22882, ZN => n4114);
   U14006 : OAI22_X1 port map( A1 => n16620, A2 => n23624, B1 => n19983, B2 => 
                           n22882, ZN => n4115);
   U14007 : OAI22_X1 port map( A1 => n16619, A2 => n23623, B1 => n19982, B2 => 
                           n22882, ZN => n4116);
   U14008 : OAI22_X1 port map( A1 => n16618, A2 => n23622, B1 => n19981, B2 => 
                           n22882, ZN => n4117);
   U14009 : OAI22_X1 port map( A1 => n16617, A2 => n23624, B1 => n19980, B2 => 
                           n22882, ZN => n4118);
   U14010 : OAI22_X1 port map( A1 => n16611, A2 => n23622, B1 => n19974, B2 => 
                           n22883, ZN => n4124);
   U14011 : OAI22_X1 port map( A1 => n16610, A2 => n23622, B1 => n19973, B2 => 
                           n22883, ZN => n4125);
   U14012 : OAI22_X1 port map( A1 => n16609, A2 => n23624, B1 => n19972, B2 => 
                           n22883, ZN => n4126);
   U14013 : OAI22_X1 port map( A1 => n16608, A2 => n23623, B1 => n19971, B2 => 
                           n22883, ZN => n4127);
   U14014 : OAI22_X1 port map( A1 => n16607, A2 => n23622, B1 => n19970, B2 => 
                           n22883, ZN => n4128);
   U14015 : OAI22_X1 port map( A1 => n16606, A2 => n23622, B1 => n19969, B2 => 
                           n22883, ZN => n4129);
   U14016 : OAI22_X1 port map( A1 => n16605, A2 => n23624, B1 => n19968, B2 => 
                           n22883, ZN => n4130);
   U14017 : OAI22_X1 port map( A1 => n16635, A2 => n23642, B1 => n19870, B2 => 
                           n22893, ZN => n4228);
   U14018 : OAI22_X1 port map( A1 => n16634, A2 => n23642, B1 => n19869, B2 => 
                           n22893, ZN => n4229);
   U14019 : OAI22_X1 port map( A1 => n16633, A2 => n23642, B1 => n19868, B2 => 
                           n22893, ZN => n4230);
   U14020 : OAI22_X1 port map( A1 => n16632, A2 => n23642, B1 => n19867, B2 => 
                           n22893, ZN => n4231);
   U14021 : OAI22_X1 port map( A1 => n16631, A2 => n23642, B1 => n19866, B2 => 
                           n22893, ZN => n4232);
   U14022 : OAI22_X1 port map( A1 => n16630, A2 => n23642, B1 => n19865, B2 => 
                           n22893, ZN => n4233);
   U14023 : OAI22_X1 port map( A1 => n16629, A2 => n23642, B1 => n19864, B2 => 
                           n22893, ZN => n4234);
   U14024 : OAI22_X1 port map( A1 => n16623, A2 => n23644, B1 => n19858, B2 => 
                           n22894, ZN => n4240);
   U14025 : OAI22_X1 port map( A1 => n16622, A2 => n23643, B1 => n19857, B2 => 
                           n22894, ZN => n4241);
   U14026 : OAI22_X1 port map( A1 => n16621, A2 => n23642, B1 => n19856, B2 => 
                           n22894, ZN => n4242);
   U14027 : OAI22_X1 port map( A1 => n16620, A2 => n23644, B1 => n19855, B2 => 
                           n22894, ZN => n4243);
   U14028 : OAI22_X1 port map( A1 => n16619, A2 => n23643, B1 => n19854, B2 => 
                           n22894, ZN => n4244);
   U14029 : OAI22_X1 port map( A1 => n16618, A2 => n23642, B1 => n19853, B2 => 
                           n22894, ZN => n4245);
   U14030 : OAI22_X1 port map( A1 => n16617, A2 => n23644, B1 => n19852, B2 => 
                           n22894, ZN => n4246);
   U14031 : OAI22_X1 port map( A1 => n16611, A2 => n23642, B1 => n19846, B2 => 
                           n22895, ZN => n4252);
   U14032 : OAI22_X1 port map( A1 => n16610, A2 => n23642, B1 => n19845, B2 => 
                           n22895, ZN => n4253);
   U14033 : OAI22_X1 port map( A1 => n16609, A2 => n23644, B1 => n19844, B2 => 
                           n22895, ZN => n4254);
   U14034 : OAI22_X1 port map( A1 => n16608, A2 => n23643, B1 => n19843, B2 => 
                           n22895, ZN => n4255);
   U14035 : OAI22_X1 port map( A1 => n16607, A2 => n23642, B1 => n19842, B2 => 
                           n22895, ZN => n4256);
   U14036 : OAI22_X1 port map( A1 => n16606, A2 => n23642, B1 => n19841, B2 => 
                           n22895, ZN => n4257);
   U14037 : OAI22_X1 port map( A1 => n16605, A2 => n23644, B1 => n19840, B2 => 
                           n22895, ZN => n4258);
   U14038 : OAI22_X1 port map( A1 => n16635, A2 => n23662, B1 => n19742, B2 => 
                           n22905, ZN => n4356);
   U14039 : OAI22_X1 port map( A1 => n16634, A2 => n23662, B1 => n19741, B2 => 
                           n22905, ZN => n4357);
   U14040 : OAI22_X1 port map( A1 => n16633, A2 => n23662, B1 => n19740, B2 => 
                           n22905, ZN => n4358);
   U14041 : OAI22_X1 port map( A1 => n16632, A2 => n23662, B1 => n19739, B2 => 
                           n22905, ZN => n4359);
   U14042 : OAI22_X1 port map( A1 => n16631, A2 => n23662, B1 => n19738, B2 => 
                           n22905, ZN => n4360);
   U14043 : OAI22_X1 port map( A1 => n16630, A2 => n23662, B1 => n19737, B2 => 
                           n22905, ZN => n4361);
   U14044 : OAI22_X1 port map( A1 => n16629, A2 => n23662, B1 => n19736, B2 => 
                           n22905, ZN => n4362);
   U14045 : OAI22_X1 port map( A1 => n16623, A2 => n23664, B1 => n19730, B2 => 
                           n22906, ZN => n4368);
   U14046 : OAI22_X1 port map( A1 => n16622, A2 => n23663, B1 => n19729, B2 => 
                           n22906, ZN => n4369);
   U14047 : OAI22_X1 port map( A1 => n16621, A2 => n23662, B1 => n19728, B2 => 
                           n22906, ZN => n4370);
   U14048 : OAI22_X1 port map( A1 => n16620, A2 => n23664, B1 => n19727, B2 => 
                           n22906, ZN => n4371);
   U14049 : OAI22_X1 port map( A1 => n16619, A2 => n23663, B1 => n19726, B2 => 
                           n22906, ZN => n4372);
   U14050 : OAI22_X1 port map( A1 => n16618, A2 => n23662, B1 => n19725, B2 => 
                           n22906, ZN => n4373);
   U14051 : OAI22_X1 port map( A1 => n16617, A2 => n23664, B1 => n19724, B2 => 
                           n22906, ZN => n4374);
   U14052 : OAI22_X1 port map( A1 => n16611, A2 => n23662, B1 => n19718, B2 => 
                           n22907, ZN => n4380);
   U14053 : OAI22_X1 port map( A1 => n16610, A2 => n23662, B1 => n19717, B2 => 
                           n22907, ZN => n4381);
   U14054 : OAI22_X1 port map( A1 => n16609, A2 => n23664, B1 => n19716, B2 => 
                           n22907, ZN => n4382);
   U14055 : OAI22_X1 port map( A1 => n16608, A2 => n23663, B1 => n19715, B2 => 
                           n22907, ZN => n4383);
   U14056 : OAI22_X1 port map( A1 => n16607, A2 => n23662, B1 => n19714, B2 => 
                           n22907, ZN => n4384);
   U14057 : OAI22_X1 port map( A1 => n16606, A2 => n23662, B1 => n19713, B2 => 
                           n22907, ZN => n4385);
   U14058 : OAI22_X1 port map( A1 => n16605, A2 => n23664, B1 => n19712, B2 => 
                           n22907, ZN => n4386);
   U14059 : AOI221_X1 port map( B1 => n23867, B2 => n21259, C1 => n23851, C2 =>
                           n21743, A => n16287, ZN => n16286);
   U14060 : OAI22_X1 port map( A1 => n18998, A2 => n23311, B1 => n19126, B2 => 
                           n23325, ZN => n16287);
   U14061 : AOI221_X1 port map( B1 => n23867, B2 => n21258, C1 => n23851, C2 =>
                           n21742, A => n16266, ZN => n16265);
   U14062 : OAI22_X1 port map( A1 => n18946, A2 => n23311, B1 => n19074, B2 => 
                           n23324, ZN => n16266);
   U14063 : AOI221_X1 port map( B1 => n23867, B2 => n21221, C1 => n23851, C2 =>
                           n21706, A => n16245, ZN => n16244);
   U14064 : OAI22_X1 port map( A1 => n18997, A2 => n23311, B1 => n19125, B2 => 
                           n23323, ZN => n16245);
   U14065 : AOI221_X1 port map( B1 => n23867, B2 => n21241, C1 => n23851, C2 =>
                           n21726, A => n16224, ZN => n16223);
   U14066 : OAI22_X1 port map( A1 => n18947, A2 => n23311, B1 => n19075, B2 => 
                           n23321, ZN => n16224);
   U14067 : AOI221_X1 port map( B1 => n23867, B2 => n21257, C1 => n23851, C2 =>
                           n21741, A => n16203, ZN => n16202);
   U14068 : OAI22_X1 port map( A1 => n18996, A2 => n23311, B1 => n19124, B2 => 
                           n23321, ZN => n16203);
   U14069 : AOI221_X1 port map( B1 => n23867, B2 => n21220, C1 => n23851, C2 =>
                           n21705, A => n16182, ZN => n16181);
   U14070 : OAI22_X1 port map( A1 => n18948, A2 => n23311, B1 => n19076, B2 => 
                           n23322, ZN => n16182);
   U14071 : AOI221_X1 port map( B1 => n23867, B2 => n21256, C1 => n23851, C2 =>
                           n21740, A => n16161, ZN => n16160);
   U14072 : OAI22_X1 port map( A1 => n18995, A2 => n23314, B1 => n19123, B2 => 
                           n23323, ZN => n16161);
   U14073 : AOI221_X1 port map( B1 => n23868, B2 => n21255, C1 => n23852, C2 =>
                           n21739, A => n16140, ZN => n16139);
   U14074 : OAI22_X1 port map( A1 => n18949, A2 => n23312, B1 => n19077, B2 => 
                           n23323, ZN => n16140);
   U14075 : AOI221_X1 port map( B1 => n23868, B2 => n21219, C1 => n23852, C2 =>
                           n21704, A => n16119, ZN => n16118);
   U14076 : OAI22_X1 port map( A1 => n18994, A2 => n23311, B1 => n19122, B2 => 
                           n23323, ZN => n16119);
   U14077 : AOI221_X1 port map( B1 => n23868, B2 => n21254, C1 => n23852, C2 =>
                           n21738, A => n16098, ZN => n16097);
   U14078 : OAI22_X1 port map( A1 => n18950, A2 => n23313, B1 => n19078, B2 => 
                           n23323, ZN => n16098);
   U14079 : AOI221_X1 port map( B1 => n23868, B2 => n21218, C1 => n23852, C2 =>
                           n21703, A => n16077, ZN => n16076);
   U14080 : OAI22_X1 port map( A1 => n18993, A2 => n23310, B1 => n19121, B2 => 
                           n23323, ZN => n16077);
   U14081 : AOI221_X1 port map( B1 => n23868, B2 => n21253, C1 => n23852, C2 =>
                           n21737, A => n16056, ZN => n16055);
   U14082 : OAI22_X1 port map( A1 => n18951, A2 => n23309, B1 => n19079, B2 => 
                           n23323, ZN => n16056);
   U14083 : AOI221_X1 port map( B1 => n23868, B2 => n21280, C1 => n23852, C2 =>
                           n21836, A => n16035, ZN => n16034);
   U14084 : OAI22_X1 port map( A1 => n18992, A2 => n23312, B1 => n19120, B2 => 
                           n23324, ZN => n16035);
   U14085 : AOI221_X1 port map( B1 => n23869, B2 => n21217, C1 => n23853, C2 =>
                           n21702, A => n16014, ZN => n16013);
   U14086 : OAI22_X1 port map( A1 => n18952, A2 => n23312, B1 => n19080, B2 => 
                           n23324, ZN => n16014);
   U14087 : AOI221_X1 port map( B1 => n23869, B2 => n21240, C1 => n23853, C2 =>
                           n21725, A => n15993, ZN => n15992);
   U14088 : OAI22_X1 port map( A1 => n18991, A2 => n23312, B1 => n19119, B2 => 
                           n23324, ZN => n15993);
   U14089 : AOI221_X1 port map( B1 => n23869, B2 => n21283, C1 => n23853, C2 =>
                           n21839, A => n15972, ZN => n15971);
   U14090 : OAI22_X1 port map( A1 => n18953, A2 => n23312, B1 => n19081, B2 => 
                           n23324, ZN => n15972);
   U14091 : AOI221_X1 port map( B1 => n23869, B2 => n21282, C1 => n23853, C2 =>
                           n21838, A => n15951, ZN => n15950);
   U14092 : OAI22_X1 port map( A1 => n18990, A2 => n23312, B1 => n19118, B2 => 
                           n23324, ZN => n15951);
   U14093 : AOI221_X1 port map( B1 => n23869, B2 => n21216, C1 => n23853, C2 =>
                           n21701, A => n15930, ZN => n15929);
   U14094 : OAI22_X1 port map( A1 => n18954, A2 => n23312, B1 => n19082, B2 => 
                           n23324, ZN => n15930);
   U14095 : AOI221_X1 port map( B1 => n23869, B2 => n21252, C1 => n23853, C2 =>
                           n21736, A => n15909, ZN => n15908);
   U14096 : OAI22_X1 port map( A1 => n18989, A2 => n23313, B1 => n19117, B2 => 
                           n23323, ZN => n15909);
   U14097 : AOI221_X1 port map( B1 => n23870, B2 => n21215, C1 => n23854, C2 =>
                           n21700, A => n15888, ZN => n15887);
   U14098 : OAI22_X1 port map( A1 => n18955, A2 => n23313, B1 => n19083, B2 => 
                           n23326, ZN => n15888);
   U14099 : AOI221_X1 port map( B1 => n23870, B2 => n21281, C1 => n23854, C2 =>
                           n21837, A => n15867, ZN => n15866);
   U14100 : OAI22_X1 port map( A1 => n18988, A2 => n23313, B1 => n19116, B2 => 
                           n23325, ZN => n15867);
   U14101 : AOI221_X1 port map( B1 => n23870, B2 => n21239, C1 => n23854, C2 =>
                           n21724, A => n15846, ZN => n15845);
   U14102 : OAI22_X1 port map( A1 => n18956, A2 => n23313, B1 => n19084, B2 => 
                           n23322, ZN => n15846);
   U14103 : AOI221_X1 port map( B1 => n23870, B2 => n21238, C1 => n23854, C2 =>
                           n21723, A => n15825, ZN => n15824);
   U14104 : OAI22_X1 port map( A1 => n18987, A2 => n23313, B1 => n19115, B2 => 
                           n23321, ZN => n15825);
   U14105 : AOI221_X1 port map( B1 => n23870, B2 => n21237, C1 => n23854, C2 =>
                           n21722, A => n15804, ZN => n15803);
   U14106 : OAI22_X1 port map( A1 => n18957, A2 => n23313, B1 => n19085, B2 => 
                           n23324, ZN => n15804);
   U14107 : AOI221_X1 port map( B1 => n23870, B2 => n21251, C1 => n23854, C2 =>
                           n21735, A => n15783, ZN => n15782);
   U14108 : OAI22_X1 port map( A1 => n18986, A2 => n23309, B1 => n19114, B2 => 
                           n23325, ZN => n15783);
   U14109 : AOI221_X1 port map( B1 => n23870, B2 => n21236, C1 => n23854, C2 =>
                           n21721, A => n15762, ZN => n15761);
   U14110 : OAI22_X1 port map( A1 => n18958, A2 => n23310, B1 => n19086, B2 => 
                           n23326, ZN => n15762);
   U14111 : AOI221_X1 port map( B1 => n23871, B2 => n21214, C1 => n23855, C2 =>
                           n21699, A => n15741, ZN => n15740);
   U14112 : OAI22_X1 port map( A1 => n18985, A2 => n23314, B1 => n19113, B2 => 
                           n23325, ZN => n15741);
   U14113 : AOI221_X1 port map( B1 => n23871, B2 => n21250, C1 => n23855, C2 =>
                           n21734, A => n15720, ZN => n15719);
   U14114 : OAI22_X1 port map( A1 => n18959, A2 => n23314, B1 => n19087, B2 => 
                           n23323, ZN => n15720);
   U14115 : AOI221_X1 port map( B1 => n23871, B2 => n21213, C1 => n23855, C2 =>
                           n21698, A => n15699, ZN => n15698);
   U14116 : OAI22_X1 port map( A1 => n18984, A2 => n23311, B1 => n19112, B2 => 
                           n23323, ZN => n15699);
   U14117 : AOI221_X1 port map( B1 => n23871, B2 => n21235, C1 => n23855, C2 =>
                           n21720, A => n15678, ZN => n15677);
   U14118 : OAI22_X1 port map( A1 => n18960, A2 => n23311, B1 => n19088, B2 => 
                           n23321, ZN => n15678);
   U14119 : AOI221_X1 port map( B1 => n23871, B2 => n21274, C1 => n23855, C2 =>
                           n21765, A => n15657, ZN => n15656);
   U14120 : OAI22_X1 port map( A1 => n18983, A2 => n23313, B1 => n19111, B2 => 
                           n23324, ZN => n15657);
   U14121 : AOI221_X1 port map( B1 => n23871, B2 => n21249, C1 => n23855, C2 =>
                           n21733, A => n15636, ZN => n15635);
   U14122 : OAI22_X1 port map( A1 => n18961, A2 => n23313, B1 => n19089, B2 => 
                           n23325, ZN => n15636);
   U14123 : AOI221_X1 port map( B1 => n23872, B2 => n21234, C1 => n23856, C2 =>
                           n21719, A => n15615, ZN => n15614);
   U14124 : OAI22_X1 port map( A1 => n18982, A2 => n23312, B1 => n19110, B2 => 
                           n23326, ZN => n15615);
   U14125 : AOI221_X1 port map( B1 => n23872, B2 => n21212, C1 => n23856, C2 =>
                           n21697, A => n15594, ZN => n15593);
   U14126 : OAI22_X1 port map( A1 => n18962, A2 => n23313, B1 => n19090, B2 => 
                           n23321, ZN => n15594);
   U14127 : AOI221_X1 port map( B1 => n23872, B2 => n21233, C1 => n23856, C2 =>
                           n21718, A => n15573, ZN => n15572);
   U14128 : OAI22_X1 port map( A1 => n18981, A2 => n23313, B1 => n19109, B2 => 
                           n23322, ZN => n15573);
   U14129 : AOI221_X1 port map( B1 => n23872, B2 => n21248, C1 => n23856, C2 =>
                           n21732, A => n15552, ZN => n15551);
   U14130 : OAI22_X1 port map( A1 => n18963, A2 => n23309, B1 => n19091, B2 => 
                           n23323, ZN => n15552);
   U14131 : AOI221_X1 port map( B1 => n23835, B2 => n21814, C1 => n23824, C2 =>
                           n22176, A => n16288, ZN => n16285);
   U14132 : OAI22_X1 port map( A1 => n18806, A2 => n23288, B1 => n18934, B2 => 
                           n23302, ZN => n16288);
   U14133 : AOI221_X1 port map( B1 => n23835, B2 => n21813, C1 => n23824, C2 =>
                           n22175, A => n16267, ZN => n16264);
   U14134 : OAI22_X1 port map( A1 => n18754, A2 => n23288, B1 => n18882, B2 => 
                           n23301, ZN => n16267);
   U14135 : AOI221_X1 port map( B1 => n23835, B2 => n21812, C1 => n23824, C2 =>
                           n22174, A => n16246, ZN => n16243);
   U14136 : OAI22_X1 port map( A1 => n18805, A2 => n23288, B1 => n18933, B2 => 
                           n23300, ZN => n16246);
   U14137 : AOI221_X1 port map( B1 => n23835, B2 => n21811, C1 => n23824, C2 =>
                           n22173, A => n16225, ZN => n16222);
   U14138 : OAI22_X1 port map( A1 => n18755, A2 => n23288, B1 => n18883, B2 => 
                           n23298, ZN => n16225);
   U14139 : AOI221_X1 port map( B1 => n23835, B2 => n21810, C1 => n23823, C2 =>
                           n22054, A => n16204, ZN => n16201);
   U14140 : OAI22_X1 port map( A1 => n18804, A2 => n23288, B1 => n18932, B2 => 
                           n23298, ZN => n16204);
   U14141 : AOI221_X1 port map( B1 => n23835, B2 => n21809, C1 => n23823, C2 =>
                           n22172, A => n16183, ZN => n16180);
   U14142 : OAI22_X1 port map( A1 => n18756, A2 => n23288, B1 => n18884, B2 => 
                           n23299, ZN => n16183);
   U14143 : AOI221_X1 port map( B1 => n23835, B2 => n21808, C1 => n23823, C2 =>
                           n22171, A => n16162, ZN => n16159);
   U14144 : OAI22_X1 port map( A1 => n18803, A2 => n23291, B1 => n18931, B2 => 
                           n23300, ZN => n16162);
   U14145 : AOI221_X1 port map( B1 => n23836, B2 => n21807, C1 => n23823, C2 =>
                           n22170, A => n16141, ZN => n16138);
   U14146 : OAI22_X1 port map( A1 => n18757, A2 => n23289, B1 => n18885, B2 => 
                           n23300, ZN => n16141);
   U14147 : AOI221_X1 port map( B1 => n23836, B2 => n21806, C1 => n23823, C2 =>
                           n22169, A => n16120, ZN => n16117);
   U14148 : OAI22_X1 port map( A1 => n18802, A2 => n23288, B1 => n18930, B2 => 
                           n23300, ZN => n16120);
   U14149 : AOI221_X1 port map( B1 => n23836, B2 => n21805, C1 => n23823, C2 =>
                           n22168, A => n16099, ZN => n16096);
   U14150 : OAI22_X1 port map( A1 => n18758, A2 => n23290, B1 => n18886, B2 => 
                           n23300, ZN => n16099);
   U14151 : AOI221_X1 port map( B1 => n23836, B2 => n21804, C1 => n23822, C2 =>
                           n22167, A => n16078, ZN => n16075);
   U14152 : OAI22_X1 port map( A1 => n18801, A2 => n23286, B1 => n18929, B2 => 
                           n23300, ZN => n16078);
   U14153 : AOI221_X1 port map( B1 => n23836, B2 => n21803, C1 => n23822, C2 =>
                           n22053, A => n16057, ZN => n16054);
   U14154 : OAI22_X1 port map( A1 => n18759, A2 => n23287, B1 => n18887, B2 => 
                           n23300, ZN => n16057);
   U14155 : AOI221_X1 port map( B1 => n23836, B2 => n21802, C1 => n23822, C2 =>
                           n22166, A => n16036, ZN => n16033);
   U14156 : OAI22_X1 port map( A1 => n18800, A2 => n23289, B1 => n18928, B2 => 
                           n23301, ZN => n16036);
   U14157 : AOI221_X1 port map( B1 => n23837, B2 => n21801, C1 => n23822, C2 =>
                           n22165, A => n16015, ZN => n16012);
   U14158 : OAI22_X1 port map( A1 => n18760, A2 => n23289, B1 => n18888, B2 => 
                           n23301, ZN => n16015);
   U14159 : AOI221_X1 port map( B1 => n23837, B2 => n21800, C1 => n23822, C2 =>
                           n22052, A => n15994, ZN => n15991);
   U14160 : OAI22_X1 port map( A1 => n18799, A2 => n23289, B1 => n18927, B2 => 
                           n23301, ZN => n15994);
   U14161 : AOI221_X1 port map( B1 => n23837, B2 => n21799, C1 => n23822, C2 =>
                           n22164, A => n15973, ZN => n15970);
   U14162 : OAI22_X1 port map( A1 => n18761, A2 => n23289, B1 => n18889, B2 => 
                           n23301, ZN => n15973);
   U14163 : AOI221_X1 port map( B1 => n23837, B2 => n21798, C1 => n23821, C2 =>
                           n22163, A => n15952, ZN => n15949);
   U14164 : OAI22_X1 port map( A1 => n18798, A2 => n23289, B1 => n18926, B2 => 
                           n23301, ZN => n15952);
   U14165 : AOI221_X1 port map( B1 => n23837, B2 => n21797, C1 => n23821, C2 =>
                           n22162, A => n15931, ZN => n15928);
   U14166 : OAI22_X1 port map( A1 => n18762, A2 => n23289, B1 => n18890, B2 => 
                           n23301, ZN => n15931);
   U14167 : AOI221_X1 port map( B1 => n23837, B2 => n21796, C1 => n23821, C2 =>
                           n22161, A => n15910, ZN => n15907);
   U14168 : OAI22_X1 port map( A1 => n18797, A2 => n23290, B1 => n18925, B2 => 
                           n23300, ZN => n15910);
   U14169 : AOI221_X1 port map( B1 => n23838, B2 => n21795, C1 => n23821, C2 =>
                           n22051, A => n15889, ZN => n15886);
   U14170 : OAI22_X1 port map( A1 => n18763, A2 => n23290, B1 => n18891, B2 => 
                           n23299, ZN => n15889);
   U14171 : AOI221_X1 port map( B1 => n23838, B2 => n21794, C1 => n23821, C2 =>
                           n22050, A => n15868, ZN => n15865);
   U14172 : OAI22_X1 port map( A1 => n18796, A2 => n23290, B1 => n18924, B2 => 
                           n23303, ZN => n15868);
   U14173 : AOI221_X1 port map( B1 => n23838, B2 => n21793, C1 => n23821, C2 =>
                           n22049, A => n15847, ZN => n15844);
   U14174 : OAI22_X1 port map( A1 => n18764, A2 => n23290, B1 => n18892, B2 => 
                           n23302, ZN => n15847);
   U14175 : AOI221_X1 port map( B1 => n23838, B2 => n21792, C1 => n23820, C2 =>
                           n22048, A => n15826, ZN => n15823);
   U14176 : OAI22_X1 port map( A1 => n18795, A2 => n23290, B1 => n18923, B2 => 
                           n23298, ZN => n15826);
   U14177 : AOI221_X1 port map( B1 => n23838, B2 => n21791, C1 => n23820, C2 =>
                           n22047, A => n15805, ZN => n15802);
   U14178 : OAI22_X1 port map( A1 => n18765, A2 => n23290, B1 => n18893, B2 => 
                           n23301, ZN => n15805);
   U14179 : AOI221_X1 port map( B1 => n23838, B2 => n21790, C1 => n23820, C2 =>
                           n22046, A => n15784, ZN => n15781);
   U14180 : OAI22_X1 port map( A1 => n18794, A2 => n23286, B1 => n18922, B2 => 
                           n23302, ZN => n15784);
   U14181 : AOI221_X1 port map( B1 => n23838, B2 => n21789, C1 => n23820, C2 =>
                           n22045, A => n15763, ZN => n15760);
   U14182 : OAI22_X1 port map( A1 => n18766, A2 => n23287, B1 => n18894, B2 => 
                           n23303, ZN => n15763);
   U14183 : AOI221_X1 port map( B1 => n23839, B2 => n21788, C1 => n23820, C2 =>
                           n22044, A => n15742, ZN => n15739);
   U14184 : OAI22_X1 port map( A1 => n18793, A2 => n23291, B1 => n18921, B2 => 
                           n23302, ZN => n15742);
   U14185 : AOI221_X1 port map( B1 => n23839, B2 => n21787, C1 => n23820, C2 =>
                           n22043, A => n15721, ZN => n15718);
   U14186 : OAI22_X1 port map( A1 => n18767, A2 => n23291, B1 => n18895, B2 => 
                           n23300, ZN => n15721);
   U14187 : AOI221_X1 port map( B1 => n23839, B2 => n21786, C1 => n23819, C2 =>
                           n22160, A => n15700, ZN => n15697);
   U14188 : OAI22_X1 port map( A1 => n18792, A2 => n23288, B1 => n18920, B2 => 
                           n23300, ZN => n15700);
   U14189 : AOI221_X1 port map( B1 => n23839, B2 => n21785, C1 => n23819, C2 =>
                           n22159, A => n15679, ZN => n15676);
   U14190 : OAI22_X1 port map( A1 => n18768, A2 => n23288, B1 => n18896, B2 => 
                           n23298, ZN => n15679);
   U14191 : AOI221_X1 port map( B1 => n23839, B2 => n21784, C1 => n23819, C2 =>
                           n22042, A => n15658, ZN => n15655);
   U14192 : OAI22_X1 port map( A1 => n18791, A2 => n23290, B1 => n18919, B2 => 
                           n23301, ZN => n15658);
   U14193 : AOI221_X1 port map( B1 => n23839, B2 => n21783, C1 => n23819, C2 =>
                           n22158, A => n15637, ZN => n15634);
   U14194 : OAI22_X1 port map( A1 => n18769, A2 => n23290, B1 => n18897, B2 => 
                           n23302, ZN => n15637);
   U14195 : AOI221_X1 port map( B1 => n23840, B2 => n21782, C1 => n23819, C2 =>
                           n22157, A => n15616, ZN => n15613);
   U14196 : OAI22_X1 port map( A1 => n18790, A2 => n23289, B1 => n18918, B2 => 
                           n23303, ZN => n15616);
   U14197 : AOI221_X1 port map( B1 => n23840, B2 => n21781, C1 => n23819, C2 =>
                           n22156, A => n15595, ZN => n15592);
   U14198 : OAI22_X1 port map( A1 => n18770, A2 => n23290, B1 => n18898, B2 => 
                           n23298, ZN => n15595);
   U14199 : AOI221_X1 port map( B1 => n23840, B2 => n21780, C1 => n23818, C2 =>
                           n22041, A => n15574, ZN => n15571);
   U14200 : OAI22_X1 port map( A1 => n18789, A2 => n23290, B1 => n18917, B2 => 
                           n23299, ZN => n15574);
   U14201 : AOI221_X1 port map( B1 => n23840, B2 => n21779, C1 => n23818, C2 =>
                           n22155, A => n15553, ZN => n15550);
   U14202 : OAI22_X1 port map( A1 => n18771, A2 => n23286, B1 => n18899, B2 => 
                           n23300, ZN => n15553);
   U14203 : OAI22_X1 port map( A1 => n16636, A2 => n23642, B1 => n19871, B2 => 
                           n22893, ZN => n4227);
   U14204 : OAI22_X1 port map( A1 => n16628, A2 => n23642, B1 => n19863, B2 => 
                           n22896, ZN => n4235);
   U14205 : OAI22_X1 port map( A1 => n16627, A2 => n23642, B1 => n19862, B2 => 
                           n22894, ZN => n4236);
   U14206 : OAI22_X1 port map( A1 => n16626, A2 => n23642, B1 => n19861, B2 => 
                           n22894, ZN => n4237);
   U14207 : OAI22_X1 port map( A1 => n16625, A2 => n23642, B1 => n19860, B2 => 
                           n22894, ZN => n4238);
   U14208 : OAI22_X1 port map( A1 => n16624, A2 => n23643, B1 => n19859, B2 => 
                           n22894, ZN => n4239);
   U14209 : OAI22_X1 port map( A1 => n16616, A2 => n23642, B1 => n19851, B2 => 
                           n22894, ZN => n4247);
   U14210 : OAI22_X1 port map( A1 => n16615, A2 => n23644, B1 => n19850, B2 => 
                           n22895, ZN => n4248);
   U14211 : OAI22_X1 port map( A1 => n16614, A2 => n23643, B1 => n19849, B2 => 
                           n22895, ZN => n4249);
   U14212 : OAI22_X1 port map( A1 => n16613, A2 => n23642, B1 => n19848, B2 => 
                           n22895, ZN => n4250);
   U14213 : OAI22_X1 port map( A1 => n16612, A2 => n23643, B1 => n19847, B2 => 
                           n22895, ZN => n4251);
   U14214 : OAI22_X1 port map( A1 => n16604, A2 => n23642, B1 => n19839, B2 => 
                           n22895, ZN => n4259);
   U14215 : OAI22_X1 port map( A1 => n16603, A2 => n23644, B1 => n19838, B2 => 
                           n22896, ZN => n4260);
   U14216 : OAI22_X1 port map( A1 => n16602, A2 => n23644, B1 => n19837, B2 => 
                           n22896, ZN => n4261);
   U14217 : OAI22_X1 port map( A1 => n16601, A2 => n23643, B1 => n19836, B2 => 
                           n22896, ZN => n4262);
   U14218 : OAI22_X1 port map( A1 => n16636, A2 => n23662, B1 => n19743, B2 => 
                           n22905, ZN => n4355);
   U14219 : OAI22_X1 port map( A1 => n16628, A2 => n23662, B1 => n19735, B2 => 
                           n22908, ZN => n4363);
   U14220 : OAI22_X1 port map( A1 => n16627, A2 => n23662, B1 => n19734, B2 => 
                           n22906, ZN => n4364);
   U14221 : OAI22_X1 port map( A1 => n16626, A2 => n23662, B1 => n19733, B2 => 
                           n22906, ZN => n4365);
   U14222 : OAI22_X1 port map( A1 => n16625, A2 => n23662, B1 => n19732, B2 => 
                           n22906, ZN => n4366);
   U14223 : OAI22_X1 port map( A1 => n16624, A2 => n23663, B1 => n19731, B2 => 
                           n22906, ZN => n4367);
   U14224 : OAI22_X1 port map( A1 => n16616, A2 => n23662, B1 => n19723, B2 => 
                           n22906, ZN => n4375);
   U14225 : OAI22_X1 port map( A1 => n16615, A2 => n23664, B1 => n19722, B2 => 
                           n22907, ZN => n4376);
   U14226 : OAI22_X1 port map( A1 => n16614, A2 => n23663, B1 => n19721, B2 => 
                           n22907, ZN => n4377);
   U14227 : OAI22_X1 port map( A1 => n16613, A2 => n23662, B1 => n19720, B2 => 
                           n22907, ZN => n4378);
   U14228 : OAI22_X1 port map( A1 => n16612, A2 => n23663, B1 => n19719, B2 => 
                           n22907, ZN => n4379);
   U14229 : OAI22_X1 port map( A1 => n16604, A2 => n23662, B1 => n19711, B2 => 
                           n22907, ZN => n4387);
   U14230 : OAI22_X1 port map( A1 => n16603, A2 => n23664, B1 => n19710, B2 => 
                           n22908, ZN => n4388);
   U14231 : OAI22_X1 port map( A1 => n16602, A2 => n23664, B1 => n19709, B2 => 
                           n22908, ZN => n4389);
   U14232 : OAI22_X1 port map( A1 => n16601, A2 => n23663, B1 => n19708, B2 => 
                           n22908, ZN => n4390);
   U14233 : OAI22_X1 port map( A1 => n16636, A2 => n23602, B1 => n20127, B2 => 
                           n22869, ZN => n3971);
   U14234 : OAI22_X1 port map( A1 => n16628, A2 => n23602, B1 => n20119, B2 => 
                           n22872, ZN => n3979);
   U14235 : OAI22_X1 port map( A1 => n16627, A2 => n23602, B1 => n20118, B2 => 
                           n22870, ZN => n3980);
   U14236 : OAI22_X1 port map( A1 => n16626, A2 => n23602, B1 => n20117, B2 => 
                           n22870, ZN => n3981);
   U14237 : OAI22_X1 port map( A1 => n16625, A2 => n23602, B1 => n20116, B2 => 
                           n22870, ZN => n3982);
   U14238 : OAI22_X1 port map( A1 => n16624, A2 => n23603, B1 => n20115, B2 => 
                           n22870, ZN => n3983);
   U14239 : OAI22_X1 port map( A1 => n16616, A2 => n23602, B1 => n20107, B2 => 
                           n22870, ZN => n3991);
   U14240 : OAI22_X1 port map( A1 => n16615, A2 => n23604, B1 => n20106, B2 => 
                           n22871, ZN => n3992);
   U14241 : OAI22_X1 port map( A1 => n16614, A2 => n23603, B1 => n20105, B2 => 
                           n22871, ZN => n3993);
   U14242 : OAI22_X1 port map( A1 => n16613, A2 => n23602, B1 => n20104, B2 => 
                           n22871, ZN => n3994);
   U14243 : OAI22_X1 port map( A1 => n16612, A2 => n23603, B1 => n20103, B2 => 
                           n22871, ZN => n3995);
   U14244 : OAI22_X1 port map( A1 => n16604, A2 => n23602, B1 => n20095, B2 => 
                           n22871, ZN => n4003);
   U14245 : OAI22_X1 port map( A1 => n16603, A2 => n23604, B1 => n20094, B2 => 
                           n22872, ZN => n4004);
   U14246 : OAI22_X1 port map( A1 => n16602, A2 => n23604, B1 => n20093, B2 => 
                           n22872, ZN => n4005);
   U14247 : OAI22_X1 port map( A1 => n16601, A2 => n23603, B1 => n20092, B2 => 
                           n22872, ZN => n4006);
   U14248 : OAI22_X1 port map( A1 => n16636, A2 => n23622, B1 => n19999, B2 => 
                           n22881, ZN => n4099);
   U14249 : OAI22_X1 port map( A1 => n16628, A2 => n23622, B1 => n19991, B2 => 
                           n22884, ZN => n4107);
   U14250 : OAI22_X1 port map( A1 => n16627, A2 => n23622, B1 => n19990, B2 => 
                           n22882, ZN => n4108);
   U14251 : OAI22_X1 port map( A1 => n16626, A2 => n23622, B1 => n19989, B2 => 
                           n22882, ZN => n4109);
   U14252 : OAI22_X1 port map( A1 => n16625, A2 => n23622, B1 => n19988, B2 => 
                           n22882, ZN => n4110);
   U14253 : OAI22_X1 port map( A1 => n16624, A2 => n23623, B1 => n19987, B2 => 
                           n22882, ZN => n4111);
   U14254 : OAI22_X1 port map( A1 => n16616, A2 => n23622, B1 => n19979, B2 => 
                           n22882, ZN => n4119);
   U14255 : OAI22_X1 port map( A1 => n16615, A2 => n23624, B1 => n19978, B2 => 
                           n22883, ZN => n4120);
   U14256 : OAI22_X1 port map( A1 => n16614, A2 => n23623, B1 => n19977, B2 => 
                           n22883, ZN => n4121);
   U14257 : OAI22_X1 port map( A1 => n16613, A2 => n23622, B1 => n19976, B2 => 
                           n22883, ZN => n4122);
   U14258 : OAI22_X1 port map( A1 => n16612, A2 => n23623, B1 => n19975, B2 => 
                           n22883, ZN => n4123);
   U14259 : OAI22_X1 port map( A1 => n16604, A2 => n23622, B1 => n19967, B2 => 
                           n22883, ZN => n4131);
   U14260 : OAI22_X1 port map( A1 => n16603, A2 => n23624, B1 => n19966, B2 => 
                           n22884, ZN => n4132);
   U14261 : OAI22_X1 port map( A1 => n16602, A2 => n23624, B1 => n19965, B2 => 
                           n22884, ZN => n4133);
   U14262 : OAI22_X1 port map( A1 => n16601, A2 => n23623, B1 => n19964, B2 => 
                           n22884, ZN => n4134);
   U14263 : AOI221_X1 port map( B1 => n23835, B2 => n22411, C1 => n23824, C2 =>
                           n22368, A => n16292, ZN => n16289);
   U14264 : OAI22_X1 port map( A1 => n19318, A2 => n23288, B1 => n19446, B2 => 
                           n23301, ZN => n16292);
   U14265 : AOI221_X1 port map( B1 => n23835, B2 => n22312, C1 => n23824, C2 =>
                           n22293, A => n16271, ZN => n16268);
   U14266 : OAI22_X1 port map( A1 => n19266, A2 => n23288, B1 => n19394, B2 => 
                           n23300, ZN => n16271);
   U14267 : AOI221_X1 port map( B1 => n23835, B2 => n22409, C1 => n23824, C2 =>
                           n22366, A => n16250, ZN => n16247);
   U14268 : OAI22_X1 port map( A1 => n19317, A2 => n23288, B1 => n19445, B2 => 
                           n23300, ZN => n16250);
   U14269 : AOI221_X1 port map( B1 => n23837, B2 => n22313, C1 => n23824, C2 =>
                           n22294, A => n16229, ZN => n16226);
   U14270 : OAI22_X1 port map( A1 => n19267, A2 => n23288, B1 => n19395, B2 => 
                           n23298, ZN => n16229);
   U14271 : AOI221_X1 port map( B1 => n23835, B2 => n22335, C1 => n23823, C2 =>
                           n22310, A => n16208, ZN => n16205);
   U14272 : OAI22_X1 port map( A1 => n19316, A2 => n23288, B1 => n19444, B2 => 
                           n23299, ZN => n16208);
   U14273 : AOI221_X1 port map( B1 => n23835, B2 => n22314, C1 => n23823, C2 =>
                           n22295, A => n16187, ZN => n16184);
   U14274 : OAI22_X1 port map( A1 => n19268, A2 => n23288, B1 => n19396, B2 => 
                           n23303, ZN => n16187);
   U14275 : AOI221_X1 port map( B1 => n23835, B2 => n22334, C1 => n23823, C2 =>
                           n22309, A => n16166, ZN => n16163);
   U14276 : OAI22_X1 port map( A1 => n19315, A2 => n23290, B1 => n19443, B2 => 
                           n23300, ZN => n16166);
   U14277 : AOI221_X1 port map( B1 => n23836, B2 => n22315, C1 => n23823, C2 =>
                           n22296, A => n16145, ZN => n16142);
   U14278 : OAI22_X1 port map( A1 => n19269, A2 => n23289, B1 => n19397, B2 => 
                           n23300, ZN => n16145);
   U14279 : AOI221_X1 port map( B1 => n23836, B2 => n22333, C1 => n23823, C2 =>
                           n22308, A => n16124, ZN => n16121);
   U14280 : OAI22_X1 port map( A1 => n19314, A2 => n23288, B1 => n19442, B2 => 
                           n23300, ZN => n16124);
   U14281 : AOI221_X1 port map( B1 => n23836, B2 => n22377, C1 => n23823, C2 =>
                           n22339, A => n16103, ZN => n16100);
   U14282 : OAI22_X1 port map( A1 => n19270, A2 => n23290, B1 => n19398, B2 => 
                           n23300, ZN => n16103);
   U14283 : AOI221_X1 port map( B1 => n23836, B2 => n22332, C1 => n23822, C2 =>
                           n22307, A => n16082, ZN => n16079);
   U14284 : OAI22_X1 port map( A1 => n19313, A2 => n23286, B1 => n19441, B2 => 
                           n23300, ZN => n16082);
   U14285 : AOI221_X1 port map( B1 => n23836, B2 => n22382, C1 => n23822, C2 =>
                           n22340, A => n16061, ZN => n16058);
   U14286 : OAI22_X1 port map( A1 => n19271, A2 => n23287, B1 => n19399, B2 => 
                           n23300, ZN => n16061);
   U14287 : AOI221_X1 port map( B1 => n23836, B2 => n22331, C1 => n23822, C2 =>
                           n22347, A => n16040, ZN => n16037);
   U14288 : OAI22_X1 port map( A1 => n19312, A2 => n23289, B1 => n19440, B2 => 
                           n23301, ZN => n16040);
   U14289 : AOI221_X1 port map( B1 => n23836, B2 => n22383, C1 => n23822, C2 =>
                           n22341, A => n16019, ZN => n16016);
   U14290 : OAI22_X1 port map( A1 => n19272, A2 => n23289, B1 => n19400, B2 => 
                           n23301, ZN => n16019);
   U14291 : AOI221_X1 port map( B1 => n23837, B2 => n22408, C1 => n23822, C2 =>
                           n22365, A => n15998, ZN => n15995);
   U14292 : OAI22_X1 port map( A1 => n19311, A2 => n23289, B1 => n19439, B2 => 
                           n23301, ZN => n15998);
   U14293 : AOI221_X1 port map( B1 => n23837, B2 => n22384, C1 => n23822, C2 =>
                           n22342, A => n15977, ZN => n15974);
   U14294 : OAI22_X1 port map( A1 => n19273, A2 => n23289, B1 => n19401, B2 => 
                           n23301, ZN => n15977);
   U14295 : AOI221_X1 port map( B1 => n23837, B2 => n22407, C1 => n23821, C2 =>
                           n22381, A => n15956, ZN => n15953);
   U14296 : OAI22_X1 port map( A1 => n19310, A2 => n23289, B1 => n19438, B2 => 
                           n23301, ZN => n15956);
   U14297 : AOI221_X1 port map( B1 => n23837, B2 => n22385, C1 => n23821, C2 =>
                           n22380, A => n15935, ZN => n15932);
   U14298 : OAI22_X1 port map( A1 => n19274, A2 => n23289, B1 => n19402, B2 => 
                           n23301, ZN => n15935);
   U14299 : AOI221_X1 port map( B1 => n23837, B2 => n22406, C1 => n23821, C2 =>
                           n22364, A => n15914, ZN => n15911);
   U14300 : OAI22_X1 port map( A1 => n19309, A2 => n23290, B1 => n19437, B2 => 
                           n23299, ZN => n15914);
   U14301 : AOI221_X1 port map( B1 => n23837, B2 => n22386, C1 => n23821, C2 =>
                           n22359, A => n15893, ZN => n15890);
   U14302 : OAI22_X1 port map( A1 => n19275, A2 => n23290, B1 => n19403, B2 => 
                           n23303, ZN => n15893);
   U14303 : AOI221_X1 port map( B1 => n23838, B2 => n22405, C1 => n23821, C2 =>
                           n22363, A => n15872, ZN => n15869);
   U14304 : OAI22_X1 port map( A1 => n19308, A2 => n23290, B1 => n19436, B2 => 
                           n23302, ZN => n15872);
   U14305 : AOI221_X1 port map( B1 => n23838, B2 => n22316, C1 => n23821, C2 =>
                           n22343, A => n15851, ZN => n15848);
   U14306 : OAI22_X1 port map( A1 => n19276, A2 => n23290, B1 => n19404, B2 => 
                           n23298, ZN => n15851);
   U14307 : AOI221_X1 port map( B1 => n23838, B2 => n22404, C1 => n23820, C2 =>
                           n22400, A => n15830, ZN => n15827);
   U14308 : OAI22_X1 port map( A1 => n19307, A2 => n23290, B1 => n19435, B2 => 
                           n23301, ZN => n15830);
   U14309 : AOI221_X1 port map( B1 => n23838, B2 => n22317, C1 => n23820, C2 =>
                           n22297, A => n15809, ZN => n15806);
   U14310 : OAI22_X1 port map( A1 => n19277, A2 => n23290, B1 => n19405, B2 => 
                           n23300, ZN => n15809);
   U14311 : AOI221_X1 port map( B1 => n23838, B2 => n22403, C1 => n23820, C2 =>
                           n22362, A => n15788, ZN => n15785);
   U14312 : OAI22_X1 port map( A1 => n19306, A2 => n23289, B1 => n19434, B2 => 
                           n23299, ZN => n15788);
   U14313 : AOI221_X1 port map( B1 => n23838, B2 => n22318, C1 => n23820, C2 =>
                           n22298, A => n15767, ZN => n15764);
   U14314 : OAI22_X1 port map( A1 => n19278, A2 => n23290, B1 => n19406, B2 => 
                           n23301, ZN => n15767);
   U14315 : AOI221_X1 port map( B1 => n23839, B2 => n22396, C1 => n23820, C2 =>
                           n22361, A => n15746, ZN => n15743);
   U14316 : OAI22_X1 port map( A1 => n19305, A2 => n23286, B1 => n19433, B2 => 
                           n23302, ZN => n15746);
   U14317 : AOI221_X1 port map( B1 => n23839, B2 => n22319, C1 => n23820, C2 =>
                           n22299, A => n15725, ZN => n15722);
   U14318 : OAI22_X1 port map( A1 => n19279, A2 => n23287, B1 => n19407, B2 => 
                           n23300, ZN => n15725);
   U14319 : AOI221_X1 port map( B1 => n23839, B2 => n22330, C1 => n23819, C2 =>
                           n22346, A => n15704, ZN => n15701);
   U14320 : OAI22_X1 port map( A1 => n19304, A2 => n23289, B1 => n19432, B2 => 
                           n23303, ZN => n15704);
   U14321 : AOI221_X1 port map( B1 => n23839, B2 => n22320, C1 => n23819, C2 =>
                           n22300, A => n15683, ZN => n15680);
   U14322 : OAI22_X1 port map( A1 => n19280, A2 => n23288, B1 => n19408, B2 => 
                           n23302, ZN => n15683);
   U14323 : AOI221_X1 port map( B1 => n23839, B2 => n22483, C1 => n23819, C2 =>
                           n22482, A => n15662, ZN => n15659);
   U14324 : OAI22_X1 port map( A1 => n19303, A2 => n23287, B1 => n19431, B2 => 
                           n23299, ZN => n15662);
   U14325 : AOI221_X1 port map( B1 => n23839, B2 => n22378, C1 => n23819, C2 =>
                           n22344, A => n15641, ZN => n15638);
   U14326 : OAI22_X1 port map( A1 => n19281, A2 => n23288, B1 => n19409, B2 => 
                           n23301, ZN => n15641);
   U14327 : AOI221_X1 port map( B1 => n23839, B2 => n22329, C1 => n23819, C2 =>
                           n22306, A => n15620, ZN => n15617);
   U14328 : OAI22_X1 port map( A1 => n19302, A2 => n23291, B1 => n19430, B2 => 
                           n23303, ZN => n15620);
   U14329 : AOI221_X1 port map( B1 => n23840, B2 => n22321, C1 => n23819, C2 =>
                           n22398, A => n15599, ZN => n15596);
   U14330 : OAI22_X1 port map( A1 => n19282, A2 => n23289, B1 => n19410, B2 => 
                           n23298, ZN => n15599);
   U14331 : AOI221_X1 port map( B1 => n23840, B2 => n22328, C1 => n23818, C2 =>
                           n22305, A => n15578, ZN => n15575);
   U14332 : OAI22_X1 port map( A1 => n19301, A2 => n23289, B1 => n19429, B2 => 
                           n23301, ZN => n15578);
   U14333 : AOI221_X1 port map( B1 => n23840, B2 => n22387, C1 => n23818, C2 =>
                           n22399, A => n15557, ZN => n15554);
   U14334 : OAI22_X1 port map( A1 => n19283, A2 => n23291, B1 => n19411, B2 => 
                           n23299, ZN => n15557);
   U14335 : AOI221_X1 port map( B1 => n23867, B2 => n21199, C1 => n23851, C2 =>
                           n21626, A => n16291, ZN => n16290);
   U14336 : OAI22_X1 port map( A1 => n19510, A2 => n23311, B1 => n19638, B2 => 
                           n23324, ZN => n16291);
   U14337 : AOI221_X1 port map( B1 => n23867, B2 => n21198, C1 => n23851, C2 =>
                           n21625, A => n16270, ZN => n16269);
   U14338 : OAI22_X1 port map( A1 => n19458, A2 => n23311, B1 => n19586, B2 => 
                           n23323, ZN => n16270);
   U14339 : AOI221_X1 port map( B1 => n23867, B2 => n21178, C1 => n23851, C2 =>
                           n21590, A => n16249, ZN => n16248);
   U14340 : OAI22_X1 port map( A1 => n19509, A2 => n23311, B1 => n19637, B2 => 
                           n23323, ZN => n16249);
   U14341 : AOI221_X1 port map( B1 => n23869, B2 => n21192, C1 => n23853, C2 =>
                           n21610, A => n16228, ZN => n16227);
   U14342 : OAI22_X1 port map( A1 => n19459, A2 => n23311, B1 => n19587, B2 => 
                           n23321, ZN => n16228);
   U14343 : AOI221_X1 port map( B1 => n23867, B2 => n21172, C1 => n23851, C2 =>
                           n21624, A => n16207, ZN => n16206);
   U14344 : OAI22_X1 port map( A1 => n19508, A2 => n23311, B1 => n19636, B2 => 
                           n23322, ZN => n16207);
   U14345 : AOI221_X1 port map( B1 => n23867, B2 => n21177, C1 => n23851, C2 =>
                           n21589, A => n16186, ZN => n16185);
   U14346 : OAI22_X1 port map( A1 => n19460, A2 => n23311, B1 => n19588, B2 => 
                           n23326, ZN => n16186);
   U14347 : AOI221_X1 port map( B1 => n23867, B2 => n21171, C1 => n23851, C2 =>
                           n21623, A => n16165, ZN => n16164);
   U14348 : OAI22_X1 port map( A1 => n19507, A2 => n23313, B1 => n19635, B2 => 
                           n23323, ZN => n16165);
   U14349 : AOI221_X1 port map( B1 => n23868, B2 => n21197, C1 => n23852, C2 =>
                           n21622, A => n16144, ZN => n16143);
   U14350 : OAI22_X1 port map( A1 => n19461, A2 => n23312, B1 => n19589, B2 => 
                           n23323, ZN => n16144);
   U14351 : AOI221_X1 port map( B1 => n23868, B2 => n21157, C1 => n23852, C2 =>
                           n21588, A => n16123, ZN => n16122);
   U14352 : OAI22_X1 port map( A1 => n19506, A2 => n23311, B1 => n19634, B2 => 
                           n23323, ZN => n16123);
   U14353 : AOI221_X1 port map( B1 => n23868, B2 => n21170, C1 => n23852, C2 =>
                           n21621, A => n16102, ZN => n16101);
   U14354 : OAI22_X1 port map( A1 => n19462, A2 => n23313, B1 => n19590, B2 => 
                           n23323, ZN => n16102);
   U14355 : AOI221_X1 port map( B1 => n23868, B2 => n21156, C1 => n23852, C2 =>
                           n21587, A => n16081, ZN => n16080);
   U14356 : OAI22_X1 port map( A1 => n19505, A2 => n23310, B1 => n19633, B2 => 
                           n23323, ZN => n16081);
   U14357 : AOI221_X1 port map( B1 => n23868, B2 => n21169, C1 => n23852, C2 =>
                           n21620, A => n16060, ZN => n16059);
   U14358 : OAI22_X1 port map( A1 => n19463, A2 => n23309, B1 => n19591, B2 => 
                           n23323, ZN => n16060);
   U14359 : AOI221_X1 port map( B1 => n23868, B2 => n21273, C1 => n23852, C2 =>
                           n21759, A => n16039, ZN => n16038);
   U14360 : OAI22_X1 port map( A1 => n19504, A2 => n23312, B1 => n19632, B2 => 
                           n23324, ZN => n16039);
   U14361 : AOI221_X1 port map( B1 => n23868, B2 => n21155, C1 => n23852, C2 =>
                           n21586, A => n16018, ZN => n16017);
   U14362 : OAI22_X1 port map( A1 => n19464, A2 => n23312, B1 => n19592, B2 => 
                           n23324, ZN => n16018);
   U14363 : AOI221_X1 port map( B1 => n23869, B2 => n21191, C1 => n23853, C2 =>
                           n21609, A => n15997, ZN => n15996);
   U14364 : OAI22_X1 port map( A1 => n19503, A2 => n23312, B1 => n19631, B2 => 
                           n23324, ZN => n15997);
   U14365 : AOI221_X1 port map( B1 => n23869, B2 => n21277, C1 => n23853, C2 =>
                           n21762, A => n15976, ZN => n15975);
   U14366 : OAI22_X1 port map( A1 => n19465, A2 => n23312, B1 => n19593, B2 => 
                           n23324, ZN => n15976);
   U14367 : AOI221_X1 port map( B1 => n23869, B2 => n21276, C1 => n23853, C2 =>
                           n21761, A => n15955, ZN => n15954);
   U14368 : OAI22_X1 port map( A1 => n19502, A2 => n23312, B1 => n19630, B2 => 
                           n23324, ZN => n15955);
   U14369 : AOI221_X1 port map( B1 => n23869, B2 => n21154, C1 => n23853, C2 =>
                           n21585, A => n15934, ZN => n15933);
   U14370 : OAI22_X1 port map( A1 => n19466, A2 => n23312, B1 => n19594, B2 => 
                           n23324, ZN => n15934);
   U14371 : AOI221_X1 port map( B1 => n23869, B2 => n21168, C1 => n23853, C2 =>
                           n21619, A => n15913, ZN => n15912);
   U14372 : OAI22_X1 port map( A1 => n19501, A2 => n23313, B1 => n19629, B2 => 
                           n23326, ZN => n15913);
   U14373 : AOI221_X1 port map( B1 => n23869, B2 => n21153, C1 => n23853, C2 =>
                           n21584, A => n15892, ZN => n15891);
   U14374 : OAI22_X1 port map( A1 => n19467, A2 => n23313, B1 => n19595, B2 => 
                           n23325, ZN => n15892);
   U14375 : AOI221_X1 port map( B1 => n23870, B2 => n21275, C1 => n23854, C2 =>
                           n21760, A => n15871, ZN => n15870);
   U14376 : OAI22_X1 port map( A1 => n19500, A2 => n23313, B1 => n19628, B2 => 
                           n23322, ZN => n15871);
   U14377 : AOI221_X1 port map( B1 => n23870, B2 => n21163, C1 => n23854, C2 =>
                           n21608, A => n15850, ZN => n15849);
   U14378 : OAI22_X1 port map( A1 => n19468, A2 => n23313, B1 => n19596, B2 => 
                           n23321, ZN => n15850);
   U14379 : AOI221_X1 port map( B1 => n23870, B2 => n21190, C1 => n23854, C2 =>
                           n21607, A => n15829, ZN => n15828);
   U14380 : OAI22_X1 port map( A1 => n19499, A2 => n23313, B1 => n19627, B2 => 
                           n23324, ZN => n15829);
   U14381 : AOI221_X1 port map( B1 => n23870, B2 => n21189, C1 => n23854, C2 =>
                           n21606, A => n15808, ZN => n15807);
   U14382 : OAI22_X1 port map( A1 => n19469, A2 => n23313, B1 => n19597, B2 => 
                           n23323, ZN => n15808);
   U14383 : AOI221_X1 port map( B1 => n23870, B2 => n21196, C1 => n23854, C2 =>
                           n21618, A => n15787, ZN => n15786);
   U14384 : OAI22_X1 port map( A1 => n19498, A2 => n23312, B1 => n19626, B2 => 
                           n23322, ZN => n15787);
   U14385 : AOI221_X1 port map( B1 => n23870, B2 => n21162, C1 => n23854, C2 =>
                           n21605, A => n15766, ZN => n15765);
   U14386 : OAI22_X1 port map( A1 => n19470, A2 => n23313, B1 => n19598, B2 => 
                           n23324, ZN => n15766);
   U14387 : AOI221_X1 port map( B1 => n23871, B2 => n21176, C1 => n23855, C2 =>
                           n21583, A => n15745, ZN => n15744);
   U14388 : OAI22_X1 port map( A1 => n19497, A2 => n23312, B1 => n19625, B2 => 
                           n23325, ZN => n15745);
   U14389 : AOI221_X1 port map( B1 => n23871, B2 => n21195, C1 => n23855, C2 =>
                           n21617, A => n15724, ZN => n15723);
   U14390 : OAI22_X1 port map( A1 => n19471, A2 => n23309, B1 => n19599, B2 => 
                           n23323, ZN => n15724);
   U14391 : AOI221_X1 port map( B1 => n23871, B2 => n21175, C1 => n23855, C2 =>
                           n21582, A => n15703, ZN => n15702);
   U14392 : OAI22_X1 port map( A1 => n19496, A2 => n23310, B1 => n19624, B2 => 
                           n23326, ZN => n15703);
   U14393 : AOI221_X1 port map( B1 => n23871, B2 => n21161, C1 => n23855, C2 =>
                           n21604, A => n15682, ZN => n15681);
   U14394 : OAI22_X1 port map( A1 => n19472, A2 => n23311, B1 => n19600, B2 => 
                           n23325, ZN => n15682);
   U14395 : AOI221_X1 port map( B1 => n23871, B2 => n21209, C1 => n23855, C2 =>
                           n21638, A => n15661, ZN => n15660);
   U14396 : OAI22_X1 port map( A1 => n19495, A2 => n23310, B1 => n19623, B2 => 
                           n23321, ZN => n15661);
   U14397 : AOI221_X1 port map( B1 => n23871, B2 => n21167, C1 => n23855, C2 =>
                           n21616, A => n15640, ZN => n15639);
   U14398 : OAI22_X1 port map( A1 => n19473, A2 => n23311, B1 => n19601, B2 => 
                           n23322, ZN => n15640);
   U14399 : AOI221_X1 port map( B1 => n23871, B2 => n21188, C1 => n23855, C2 =>
                           n21603, A => n15619, ZN => n15618);
   U14400 : OAI22_X1 port map( A1 => n19494, A2 => n23314, B1 => n19622, B2 => 
                           n23326, ZN => n15619);
   U14401 : AOI221_X1 port map( B1 => n23872, B2 => n21152, C1 => n23856, C2 =>
                           n21581, A => n15598, ZN => n15597);
   U14402 : OAI22_X1 port map( A1 => n19474, A2 => n23312, B1 => n19602, B2 => 
                           n23324, ZN => n15598);
   U14403 : AOI221_X1 port map( B1 => n23872, B2 => n21160, C1 => n23856, C2 =>
                           n21602, A => n15577, ZN => n15576);
   U14404 : OAI22_X1 port map( A1 => n19493, A2 => n23312, B1 => n19621, B2 => 
                           n23324, ZN => n15577);
   U14405 : AOI221_X1 port map( B1 => n23872, B2 => n21166, C1 => n23856, C2 =>
                           n21615, A => n15556, ZN => n15555);
   U14406 : OAI22_X1 port map( A1 => n19475, A2 => n23314, B1 => n19603, B2 => 
                           n23322, ZN => n15556);
   U14407 : OAI22_X1 port map( A1 => n16635, A2 => n23652, B1 => n19806, B2 => 
                           n22899, ZN => n4292);
   U14408 : OAI22_X1 port map( A1 => n16634, A2 => n23652, B1 => n19805, B2 => 
                           n22899, ZN => n4293);
   U14409 : OAI22_X1 port map( A1 => n16633, A2 => n23652, B1 => n19804, B2 => 
                           n22899, ZN => n4294);
   U14410 : OAI22_X1 port map( A1 => n16632, A2 => n23652, B1 => n19803, B2 => 
                           n22899, ZN => n4295);
   U14411 : OAI22_X1 port map( A1 => n16631, A2 => n23652, B1 => n19802, B2 => 
                           n22899, ZN => n4296);
   U14412 : OAI22_X1 port map( A1 => n16630, A2 => n23652, B1 => n19801, B2 => 
                           n22899, ZN => n4297);
   U14413 : OAI22_X1 port map( A1 => n16629, A2 => n23652, B1 => n19800, B2 => 
                           n22899, ZN => n4298);
   U14414 : OAI22_X1 port map( A1 => n16623, A2 => n23654, B1 => n19794, B2 => 
                           n22900, ZN => n4304);
   U14415 : OAI22_X1 port map( A1 => n16622, A2 => n23653, B1 => n19793, B2 => 
                           n22900, ZN => n4305);
   U14416 : OAI22_X1 port map( A1 => n16621, A2 => n23652, B1 => n19792, B2 => 
                           n22900, ZN => n4306);
   U14417 : OAI22_X1 port map( A1 => n16620, A2 => n23654, B1 => n19791, B2 => 
                           n22900, ZN => n4307);
   U14418 : OAI22_X1 port map( A1 => n16619, A2 => n23653, B1 => n19790, B2 => 
                           n22900, ZN => n4308);
   U14419 : OAI22_X1 port map( A1 => n16618, A2 => n23652, B1 => n19789, B2 => 
                           n22900, ZN => n4309);
   U14420 : OAI22_X1 port map( A1 => n16617, A2 => n23654, B1 => n19788, B2 => 
                           n22900, ZN => n4310);
   U14421 : OAI22_X1 port map( A1 => n16611, A2 => n23652, B1 => n19782, B2 => 
                           n22901, ZN => n4316);
   U14422 : OAI22_X1 port map( A1 => n16610, A2 => n23652, B1 => n19781, B2 => 
                           n22901, ZN => n4317);
   U14423 : OAI22_X1 port map( A1 => n16609, A2 => n23654, B1 => n19780, B2 => 
                           n22901, ZN => n4318);
   U14424 : OAI22_X1 port map( A1 => n16608, A2 => n23653, B1 => n19779, B2 => 
                           n22901, ZN => n4319);
   U14425 : OAI22_X1 port map( A1 => n16607, A2 => n23652, B1 => n19778, B2 => 
                           n22901, ZN => n4320);
   U14426 : OAI22_X1 port map( A1 => n16606, A2 => n23652, B1 => n19777, B2 => 
                           n22901, ZN => n4321);
   U14427 : OAI22_X1 port map( A1 => n16605, A2 => n23654, B1 => n19776, B2 => 
                           n22901, ZN => n4322);
   U14428 : OAI22_X1 port map( A1 => n16636, A2 => n23652, B1 => n19807, B2 => 
                           n22899, ZN => n4291);
   U14429 : OAI22_X1 port map( A1 => n16628, A2 => n23652, B1 => n19799, B2 => 
                           n22902, ZN => n4299);
   U14430 : OAI22_X1 port map( A1 => n16627, A2 => n23652, B1 => n19798, B2 => 
                           n22900, ZN => n4300);
   U14431 : OAI22_X1 port map( A1 => n16626, A2 => n23652, B1 => n19797, B2 => 
                           n22900, ZN => n4301);
   U14432 : OAI22_X1 port map( A1 => n16625, A2 => n23652, B1 => n19796, B2 => 
                           n22900, ZN => n4302);
   U14433 : OAI22_X1 port map( A1 => n16624, A2 => n23653, B1 => n19795, B2 => 
                           n22900, ZN => n4303);
   U14434 : OAI22_X1 port map( A1 => n16616, A2 => n23652, B1 => n19787, B2 => 
                           n22900, ZN => n4311);
   U14435 : OAI22_X1 port map( A1 => n16615, A2 => n23654, B1 => n19786, B2 => 
                           n22901, ZN => n4312);
   U14436 : OAI22_X1 port map( A1 => n16614, A2 => n23653, B1 => n19785, B2 => 
                           n22901, ZN => n4313);
   U14437 : OAI22_X1 port map( A1 => n16613, A2 => n23652, B1 => n19784, B2 => 
                           n22901, ZN => n4314);
   U14438 : OAI22_X1 port map( A1 => n16612, A2 => n23653, B1 => n19783, B2 => 
                           n22901, ZN => n4315);
   U14439 : OAI22_X1 port map( A1 => n16604, A2 => n23652, B1 => n19775, B2 => 
                           n22901, ZN => n4323);
   U14440 : OAI22_X1 port map( A1 => n16603, A2 => n23654, B1 => n19774, B2 => 
                           n22902, ZN => n4324);
   U14441 : OAI22_X1 port map( A1 => n16602, A2 => n23654, B1 => n19773, B2 => 
                           n22902, ZN => n4325);
   U14442 : OAI22_X1 port map( A1 => n16601, A2 => n23653, B1 => n19772, B2 => 
                           n22902, ZN => n4326);
   U14443 : OAI22_X1 port map( A1 => n16658, A2 => n23524, B1 => n20661, B2 => 
                           n22819, ZN => n3437);
   U14444 : OAI22_X1 port map( A1 => n16657, A2 => n23524, B1 => n20660, B2 => 
                           n22819, ZN => n3438);
   U14445 : OAI22_X1 port map( A1 => n16656, A2 => n23524, B1 => n20659, B2 => 
                           n22819, ZN => n3439);
   U14446 : OAI22_X1 port map( A1 => n16655, A2 => n23524, B1 => n20658, B2 => 
                           n22819, ZN => n3440);
   U14447 : OAI22_X1 port map( A1 => n16654, A2 => n23524, B1 => n20657, B2 => 
                           n22819, ZN => n3441);
   U14448 : OAI22_X1 port map( A1 => n16653, A2 => n23524, B1 => n20656, B2 => 
                           n22819, ZN => n3442);
   U14449 : OAI22_X1 port map( A1 => n16652, A2 => n23524, B1 => n20655, B2 => 
                           n22820, ZN => n3443);
   U14450 : OAI22_X1 port map( A1 => n16646, A2 => n23523, B1 => n20649, B2 => 
                           n22820, ZN => n3449);
   U14451 : OAI22_X1 port map( A1 => n16645, A2 => n23523, B1 => n20648, B2 => 
                           n22820, ZN => n3450);
   U14452 : OAI22_X1 port map( A1 => n16644, A2 => n23523, B1 => n20647, B2 => 
                           n22820, ZN => n3451);
   U14453 : OAI22_X1 port map( A1 => n16643, A2 => n23523, B1 => n20646, B2 => 
                           n22820, ZN => n3452);
   U14454 : OAI22_X1 port map( A1 => n16642, A2 => n23523, B1 => n20645, B2 => 
                           n22820, ZN => n3453);
   U14455 : OAI22_X1 port map( A1 => n16641, A2 => n23523, B1 => n20644, B2 => 
                           n22820, ZN => n3454);
   U14456 : OAI22_X1 port map( A1 => n16640, A2 => n23523, B1 => n20643, B2 => 
                           n22821, ZN => n3455);
   U14457 : OAI22_X1 port map( A1 => n16658, A2 => n23544, B1 => n20533, B2 => 
                           n22831, ZN => n3565);
   U14458 : OAI22_X1 port map( A1 => n16657, A2 => n23544, B1 => n20532, B2 => 
                           n22831, ZN => n3566);
   U14459 : OAI22_X1 port map( A1 => n16656, A2 => n23544, B1 => n20531, B2 => 
                           n22831, ZN => n3567);
   U14460 : OAI22_X1 port map( A1 => n16655, A2 => n23544, B1 => n20530, B2 => 
                           n22831, ZN => n3568);
   U14461 : OAI22_X1 port map( A1 => n16654, A2 => n23544, B1 => n20529, B2 => 
                           n22831, ZN => n3569);
   U14462 : OAI22_X1 port map( A1 => n16653, A2 => n23544, B1 => n20528, B2 => 
                           n22831, ZN => n3570);
   U14463 : OAI22_X1 port map( A1 => n16652, A2 => n23544, B1 => n20527, B2 => 
                           n22832, ZN => n3571);
   U14464 : OAI22_X1 port map( A1 => n16646, A2 => n23543, B1 => n20521, B2 => 
                           n22832, ZN => n3577);
   U14465 : OAI22_X1 port map( A1 => n16645, A2 => n23543, B1 => n20520, B2 => 
                           n22832, ZN => n3578);
   U14466 : OAI22_X1 port map( A1 => n16644, A2 => n23543, B1 => n20519, B2 => 
                           n22832, ZN => n3579);
   U14467 : OAI22_X1 port map( A1 => n16643, A2 => n23543, B1 => n20518, B2 => 
                           n22832, ZN => n3580);
   U14468 : OAI22_X1 port map( A1 => n16642, A2 => n23543, B1 => n20517, B2 => 
                           n22832, ZN => n3581);
   U14469 : OAI22_X1 port map( A1 => n16641, A2 => n23543, B1 => n20516, B2 => 
                           n22832, ZN => n3582);
   U14470 : OAI22_X1 port map( A1 => n16640, A2 => n23543, B1 => n20515, B2 => 
                           n22833, ZN => n3583);
   U14471 : OAI22_X1 port map( A1 => n16658, A2 => n23564, B1 => n20405, B2 => 
                           n22843, ZN => n3693);
   U14472 : OAI22_X1 port map( A1 => n16657, A2 => n23564, B1 => n20404, B2 => 
                           n22843, ZN => n3694);
   U14473 : OAI22_X1 port map( A1 => n16656, A2 => n23564, B1 => n20403, B2 => 
                           n22843, ZN => n3695);
   U14474 : OAI22_X1 port map( A1 => n16655, A2 => n23564, B1 => n20402, B2 => 
                           n22843, ZN => n3696);
   U14475 : OAI22_X1 port map( A1 => n16654, A2 => n23564, B1 => n20401, B2 => 
                           n22843, ZN => n3697);
   U14476 : OAI22_X1 port map( A1 => n16653, A2 => n23564, B1 => n20400, B2 => 
                           n22843, ZN => n3698);
   U14477 : OAI22_X1 port map( A1 => n16652, A2 => n23564, B1 => n20399, B2 => 
                           n22844, ZN => n3699);
   U14478 : OAI22_X1 port map( A1 => n16646, A2 => n23563, B1 => n20393, B2 => 
                           n22844, ZN => n3705);
   U14479 : OAI22_X1 port map( A1 => n16645, A2 => n23563, B1 => n20392, B2 => 
                           n22844, ZN => n3706);
   U14480 : OAI22_X1 port map( A1 => n16644, A2 => n23563, B1 => n20391, B2 => 
                           n22844, ZN => n3707);
   U14481 : OAI22_X1 port map( A1 => n16643, A2 => n23563, B1 => n20390, B2 => 
                           n22844, ZN => n3708);
   U14482 : OAI22_X1 port map( A1 => n16642, A2 => n23563, B1 => n20389, B2 => 
                           n22844, ZN => n3709);
   U14483 : OAI22_X1 port map( A1 => n16641, A2 => n23563, B1 => n20388, B2 => 
                           n22844, ZN => n3710);
   U14484 : OAI22_X1 port map( A1 => n16640, A2 => n23563, B1 => n20387, B2 => 
                           n22845, ZN => n3711);
   U14485 : OAI22_X1 port map( A1 => n16658, A2 => n23584, B1 => n20277, B2 => 
                           n22855, ZN => n3821);
   U14486 : OAI22_X1 port map( A1 => n16657, A2 => n23584, B1 => n20276, B2 => 
                           n22855, ZN => n3822);
   U14487 : OAI22_X1 port map( A1 => n16656, A2 => n23584, B1 => n20275, B2 => 
                           n22855, ZN => n3823);
   U14488 : OAI22_X1 port map( A1 => n16655, A2 => n23584, B1 => n20274, B2 => 
                           n22855, ZN => n3824);
   U14489 : OAI22_X1 port map( A1 => n16654, A2 => n23584, B1 => n20273, B2 => 
                           n22855, ZN => n3825);
   U14490 : OAI22_X1 port map( A1 => n16653, A2 => n23584, B1 => n20272, B2 => 
                           n22855, ZN => n3826);
   U14491 : OAI22_X1 port map( A1 => n16652, A2 => n23584, B1 => n20271, B2 => 
                           n22856, ZN => n3827);
   U14492 : OAI22_X1 port map( A1 => n16646, A2 => n23583, B1 => n20265, B2 => 
                           n22856, ZN => n3833);
   U14493 : OAI22_X1 port map( A1 => n16645, A2 => n23583, B1 => n20264, B2 => 
                           n22856, ZN => n3834);
   U14494 : OAI22_X1 port map( A1 => n16644, A2 => n23583, B1 => n20263, B2 => 
                           n22856, ZN => n3835);
   U14495 : OAI22_X1 port map( A1 => n16643, A2 => n23583, B1 => n20262, B2 => 
                           n22856, ZN => n3836);
   U14496 : OAI22_X1 port map( A1 => n16642, A2 => n23583, B1 => n20261, B2 => 
                           n22856, ZN => n3837);
   U14497 : OAI22_X1 port map( A1 => n16641, A2 => n23583, B1 => n20260, B2 => 
                           n22856, ZN => n3838);
   U14498 : OAI22_X1 port map( A1 => n16640, A2 => n23583, B1 => n20259, B2 => 
                           n22857, ZN => n3839);
   U14499 : OAI22_X1 port map( A1 => n16658, A2 => n23534, B1 => n20597, B2 => 
                           n22825, ZN => n3501);
   U14500 : OAI22_X1 port map( A1 => n16657, A2 => n23534, B1 => n20596, B2 => 
                           n22825, ZN => n3502);
   U14501 : OAI22_X1 port map( A1 => n16656, A2 => n23534, B1 => n20595, B2 => 
                           n22825, ZN => n3503);
   U14502 : OAI22_X1 port map( A1 => n16655, A2 => n23534, B1 => n20594, B2 => 
                           n22825, ZN => n3504);
   U14503 : OAI22_X1 port map( A1 => n16654, A2 => n23534, B1 => n20593, B2 => 
                           n22825, ZN => n3505);
   U14504 : OAI22_X1 port map( A1 => n16653, A2 => n23534, B1 => n20592, B2 => 
                           n22825, ZN => n3506);
   U14505 : OAI22_X1 port map( A1 => n16652, A2 => n23534, B1 => n20591, B2 => 
                           n22826, ZN => n3507);
   U14506 : OAI22_X1 port map( A1 => n16646, A2 => n23533, B1 => n20585, B2 => 
                           n22826, ZN => n3513);
   U14507 : OAI22_X1 port map( A1 => n16645, A2 => n23533, B1 => n20584, B2 => 
                           n22826, ZN => n3514);
   U14508 : OAI22_X1 port map( A1 => n16644, A2 => n23533, B1 => n20583, B2 => 
                           n22826, ZN => n3515);
   U14509 : OAI22_X1 port map( A1 => n16643, A2 => n23533, B1 => n20582, B2 => 
                           n22826, ZN => n3516);
   U14510 : OAI22_X1 port map( A1 => n16642, A2 => n23533, B1 => n20581, B2 => 
                           n22826, ZN => n3517);
   U14511 : OAI22_X1 port map( A1 => n16641, A2 => n23533, B1 => n20580, B2 => 
                           n22826, ZN => n3518);
   U14512 : OAI22_X1 port map( A1 => n16640, A2 => n23533, B1 => n20579, B2 => 
                           n22827, ZN => n3519);
   U14513 : OAI22_X1 port map( A1 => n16658, A2 => n23554, B1 => n20469, B2 => 
                           n22837, ZN => n3629);
   U14514 : OAI22_X1 port map( A1 => n16657, A2 => n23554, B1 => n20468, B2 => 
                           n22837, ZN => n3630);
   U14515 : OAI22_X1 port map( A1 => n16656, A2 => n23554, B1 => n20467, B2 => 
                           n22837, ZN => n3631);
   U14516 : OAI22_X1 port map( A1 => n16655, A2 => n23554, B1 => n20466, B2 => 
                           n22837, ZN => n3632);
   U14517 : OAI22_X1 port map( A1 => n16654, A2 => n23554, B1 => n20465, B2 => 
                           n22837, ZN => n3633);
   U14518 : OAI22_X1 port map( A1 => n16653, A2 => n23554, B1 => n20464, B2 => 
                           n22837, ZN => n3634);
   U14519 : OAI22_X1 port map( A1 => n16652, A2 => n23554, B1 => n20463, B2 => 
                           n22838, ZN => n3635);
   U14520 : OAI22_X1 port map( A1 => n16646, A2 => n23553, B1 => n20457, B2 => 
                           n22838, ZN => n3641);
   U14521 : OAI22_X1 port map( A1 => n16645, A2 => n23553, B1 => n20456, B2 => 
                           n22838, ZN => n3642);
   U14522 : OAI22_X1 port map( A1 => n16644, A2 => n23553, B1 => n20455, B2 => 
                           n22838, ZN => n3643);
   U14523 : OAI22_X1 port map( A1 => n16643, A2 => n23553, B1 => n20454, B2 => 
                           n22838, ZN => n3644);
   U14524 : OAI22_X1 port map( A1 => n16642, A2 => n23553, B1 => n20453, B2 => 
                           n22838, ZN => n3645);
   U14525 : OAI22_X1 port map( A1 => n16641, A2 => n23553, B1 => n20452, B2 => 
                           n22838, ZN => n3646);
   U14526 : OAI22_X1 port map( A1 => n16640, A2 => n23553, B1 => n20451, B2 => 
                           n22839, ZN => n3647);
   U14527 : OAI22_X1 port map( A1 => n16658, A2 => n23574, B1 => n20341, B2 => 
                           n22849, ZN => n3757);
   U14528 : OAI22_X1 port map( A1 => n16657, A2 => n23574, B1 => n20340, B2 => 
                           n22849, ZN => n3758);
   U14529 : OAI22_X1 port map( A1 => n16656, A2 => n23574, B1 => n20339, B2 => 
                           n22849, ZN => n3759);
   U14530 : OAI22_X1 port map( A1 => n16655, A2 => n23574, B1 => n20338, B2 => 
                           n22849, ZN => n3760);
   U14531 : OAI22_X1 port map( A1 => n16654, A2 => n23574, B1 => n20337, B2 => 
                           n22849, ZN => n3761);
   U14532 : OAI22_X1 port map( A1 => n16653, A2 => n23574, B1 => n20336, B2 => 
                           n22849, ZN => n3762);
   U14533 : OAI22_X1 port map( A1 => n16652, A2 => n23574, B1 => n20335, B2 => 
                           n22850, ZN => n3763);
   U14534 : OAI22_X1 port map( A1 => n16646, A2 => n23573, B1 => n20329, B2 => 
                           n22850, ZN => n3769);
   U14535 : OAI22_X1 port map( A1 => n16645, A2 => n23573, B1 => n20328, B2 => 
                           n22850, ZN => n3770);
   U14536 : OAI22_X1 port map( A1 => n16644, A2 => n23573, B1 => n20327, B2 => 
                           n22850, ZN => n3771);
   U14537 : OAI22_X1 port map( A1 => n16643, A2 => n23573, B1 => n20326, B2 => 
                           n22850, ZN => n3772);
   U14538 : OAI22_X1 port map( A1 => n16642, A2 => n23573, B1 => n20325, B2 => 
                           n22850, ZN => n3773);
   U14539 : OAI22_X1 port map( A1 => n16641, A2 => n23573, B1 => n20324, B2 => 
                           n22850, ZN => n3774);
   U14540 : OAI22_X1 port map( A1 => n16640, A2 => n23573, B1 => n20323, B2 => 
                           n22851, ZN => n3775);
   U14541 : OAI22_X1 port map( A1 => n16635, A2 => n23592, B1 => n20190, B2 => 
                           n22863, ZN => n3908);
   U14542 : OAI22_X1 port map( A1 => n16634, A2 => n23592, B1 => n20189, B2 => 
                           n22863, ZN => n3909);
   U14543 : OAI22_X1 port map( A1 => n16633, A2 => n23592, B1 => n20188, B2 => 
                           n22863, ZN => n3910);
   U14544 : OAI22_X1 port map( A1 => n16632, A2 => n23592, B1 => n20187, B2 => 
                           n22863, ZN => n3911);
   U14545 : OAI22_X1 port map( A1 => n16631, A2 => n23592, B1 => n20186, B2 => 
                           n22863, ZN => n3912);
   U14546 : OAI22_X1 port map( A1 => n16630, A2 => n23592, B1 => n20185, B2 => 
                           n22863, ZN => n3913);
   U14547 : OAI22_X1 port map( A1 => n16629, A2 => n23592, B1 => n20184, B2 => 
                           n22863, ZN => n3914);
   U14548 : OAI22_X1 port map( A1 => n16623, A2 => n23594, B1 => n20178, B2 => 
                           n22864, ZN => n3920);
   U14549 : OAI22_X1 port map( A1 => n16622, A2 => n23593, B1 => n20177, B2 => 
                           n22864, ZN => n3921);
   U14550 : OAI22_X1 port map( A1 => n16621, A2 => n23592, B1 => n20176, B2 => 
                           n22864, ZN => n3922);
   U14551 : OAI22_X1 port map( A1 => n16620, A2 => n23594, B1 => n20175, B2 => 
                           n22864, ZN => n3923);
   U14552 : OAI22_X1 port map( A1 => n16619, A2 => n23593, B1 => n20174, B2 => 
                           n22864, ZN => n3924);
   U14553 : OAI22_X1 port map( A1 => n16618, A2 => n23592, B1 => n20173, B2 => 
                           n22864, ZN => n3925);
   U14554 : OAI22_X1 port map( A1 => n16617, A2 => n23594, B1 => n20172, B2 => 
                           n22864, ZN => n3926);
   U14555 : OAI22_X1 port map( A1 => n16611, A2 => n23592, B1 => n20166, B2 => 
                           n22865, ZN => n3932);
   U14556 : OAI22_X1 port map( A1 => n16610, A2 => n23592, B1 => n20165, B2 => 
                           n22865, ZN => n3933);
   U14557 : OAI22_X1 port map( A1 => n16609, A2 => n23594, B1 => n20164, B2 => 
                           n22865, ZN => n3934);
   U14558 : OAI22_X1 port map( A1 => n16608, A2 => n23593, B1 => n20163, B2 => 
                           n22865, ZN => n3935);
   U14559 : OAI22_X1 port map( A1 => n16607, A2 => n23592, B1 => n20162, B2 => 
                           n22865, ZN => n3936);
   U14560 : OAI22_X1 port map( A1 => n16606, A2 => n23592, B1 => n20161, B2 => 
                           n22865, ZN => n3937);
   U14561 : OAI22_X1 port map( A1 => n16605, A2 => n23594, B1 => n20160, B2 => 
                           n22865, ZN => n3938);
   U14562 : OAI22_X1 port map( A1 => n16635, A2 => n23612, B1 => n20062, B2 => 
                           n22875, ZN => n4036);
   U14563 : OAI22_X1 port map( A1 => n16634, A2 => n23612, B1 => n20061, B2 => 
                           n22875, ZN => n4037);
   U14564 : OAI22_X1 port map( A1 => n16633, A2 => n23612, B1 => n20060, B2 => 
                           n22875, ZN => n4038);
   U14565 : OAI22_X1 port map( A1 => n16632, A2 => n23612, B1 => n20059, B2 => 
                           n22875, ZN => n4039);
   U14566 : OAI22_X1 port map( A1 => n16631, A2 => n23612, B1 => n20058, B2 => 
                           n22875, ZN => n4040);
   U14567 : OAI22_X1 port map( A1 => n16630, A2 => n23612, B1 => n20057, B2 => 
                           n22875, ZN => n4041);
   U14568 : OAI22_X1 port map( A1 => n16629, A2 => n23612, B1 => n20056, B2 => 
                           n22875, ZN => n4042);
   U14569 : OAI22_X1 port map( A1 => n16623, A2 => n23614, B1 => n20050, B2 => 
                           n22876, ZN => n4048);
   U14570 : OAI22_X1 port map( A1 => n16622, A2 => n23613, B1 => n20049, B2 => 
                           n22876, ZN => n4049);
   U14571 : OAI22_X1 port map( A1 => n16621, A2 => n23612, B1 => n20048, B2 => 
                           n22876, ZN => n4050);
   U14572 : OAI22_X1 port map( A1 => n16620, A2 => n23614, B1 => n20047, B2 => 
                           n22876, ZN => n4051);
   U14573 : OAI22_X1 port map( A1 => n16619, A2 => n23613, B1 => n20046, B2 => 
                           n22876, ZN => n4052);
   U14574 : OAI22_X1 port map( A1 => n16618, A2 => n23612, B1 => n20045, B2 => 
                           n22876, ZN => n4053);
   U14575 : OAI22_X1 port map( A1 => n16617, A2 => n23614, B1 => n20044, B2 => 
                           n22876, ZN => n4054);
   U14576 : OAI22_X1 port map( A1 => n16611, A2 => n23612, B1 => n20038, B2 => 
                           n22877, ZN => n4060);
   U14577 : OAI22_X1 port map( A1 => n16610, A2 => n23612, B1 => n20037, B2 => 
                           n22877, ZN => n4061);
   U14578 : OAI22_X1 port map( A1 => n16609, A2 => n23614, B1 => n20036, B2 => 
                           n22877, ZN => n4062);
   U14579 : OAI22_X1 port map( A1 => n16608, A2 => n23613, B1 => n20035, B2 => 
                           n22877, ZN => n4063);
   U14580 : OAI22_X1 port map( A1 => n16607, A2 => n23612, B1 => n20034, B2 => 
                           n22877, ZN => n4064);
   U14581 : OAI22_X1 port map( A1 => n16606, A2 => n23612, B1 => n20033, B2 => 
                           n22877, ZN => n4065);
   U14582 : OAI22_X1 port map( A1 => n16605, A2 => n23614, B1 => n20032, B2 => 
                           n22877, ZN => n4066);
   U14583 : OAI22_X1 port map( A1 => n16635, A2 => n23632, B1 => n19934, B2 => 
                           n22887, ZN => n4164);
   U14584 : OAI22_X1 port map( A1 => n16634, A2 => n23632, B1 => n19933, B2 => 
                           n22887, ZN => n4165);
   U14585 : OAI22_X1 port map( A1 => n16633, A2 => n23632, B1 => n19932, B2 => 
                           n22887, ZN => n4166);
   U14586 : OAI22_X1 port map( A1 => n16632, A2 => n23632, B1 => n19931, B2 => 
                           n22887, ZN => n4167);
   U14587 : OAI22_X1 port map( A1 => n16631, A2 => n23632, B1 => n19930, B2 => 
                           n22887, ZN => n4168);
   U14588 : OAI22_X1 port map( A1 => n16630, A2 => n23632, B1 => n19929, B2 => 
                           n22887, ZN => n4169);
   U14589 : OAI22_X1 port map( A1 => n16629, A2 => n23632, B1 => n19928, B2 => 
                           n22887, ZN => n4170);
   U14590 : OAI22_X1 port map( A1 => n16623, A2 => n23634, B1 => n19922, B2 => 
                           n22888, ZN => n4176);
   U14591 : OAI22_X1 port map( A1 => n16622, A2 => n23633, B1 => n19921, B2 => 
                           n22888, ZN => n4177);
   U14592 : OAI22_X1 port map( A1 => n16621, A2 => n23632, B1 => n19920, B2 => 
                           n22888, ZN => n4178);
   U14593 : OAI22_X1 port map( A1 => n16620, A2 => n23634, B1 => n19919, B2 => 
                           n22888, ZN => n4179);
   U14594 : OAI22_X1 port map( A1 => n16619, A2 => n23633, B1 => n19918, B2 => 
                           n22888, ZN => n4180);
   U14595 : OAI22_X1 port map( A1 => n16618, A2 => n23632, B1 => n19917, B2 => 
                           n22888, ZN => n4181);
   U14596 : OAI22_X1 port map( A1 => n16617, A2 => n23634, B1 => n19916, B2 => 
                           n22888, ZN => n4182);
   U14597 : OAI22_X1 port map( A1 => n16611, A2 => n23632, B1 => n19910, B2 => 
                           n22889, ZN => n4188);
   U14598 : OAI22_X1 port map( A1 => n16610, A2 => n23632, B1 => n19909, B2 => 
                           n22889, ZN => n4189);
   U14599 : OAI22_X1 port map( A1 => n16609, A2 => n23634, B1 => n19908, B2 => 
                           n22889, ZN => n4190);
   U14600 : OAI22_X1 port map( A1 => n16608, A2 => n23633, B1 => n19907, B2 => 
                           n22889, ZN => n4191);
   U14601 : OAI22_X1 port map( A1 => n16607, A2 => n23632, B1 => n19906, B2 => 
                           n22889, ZN => n4192);
   U14602 : OAI22_X1 port map( A1 => n16606, A2 => n23632, B1 => n19905, B2 => 
                           n22889, ZN => n4193);
   U14603 : OAI22_X1 port map( A1 => n16605, A2 => n23634, B1 => n19904, B2 => 
                           n22889, ZN => n4194);
   U14604 : OAI22_X1 port map( A1 => n16660, A2 => n23584, B1 => n20279, B2 => 
                           n22855, ZN => n3819);
   U14605 : OAI22_X1 port map( A1 => n16659, A2 => n23584, B1 => n20278, B2 => 
                           n22855, ZN => n3820);
   U14606 : OAI22_X1 port map( A1 => n16651, A2 => n23584, B1 => n20270, B2 => 
                           n22856, ZN => n3828);
   U14607 : OAI22_X1 port map( A1 => n16650, A2 => n23584, B1 => n20269, B2 => 
                           n22856, ZN => n3829);
   U14608 : OAI22_X1 port map( A1 => n16649, A2 => n23584, B1 => n20268, B2 => 
                           n22856, ZN => n3830);
   U14609 : OAI22_X1 port map( A1 => n16648, A2 => n23583, B1 => n20267, B2 => 
                           n22856, ZN => n3831);
   U14610 : OAI22_X1 port map( A1 => n16647, A2 => n23583, B1 => n20266, B2 => 
                           n22856, ZN => n3832);
   U14611 : OAI22_X1 port map( A1 => n16639, A2 => n23583, B1 => n20258, B2 => 
                           n22857, ZN => n3840);
   U14612 : OAI22_X1 port map( A1 => n16638, A2 => n23583, B1 => n20257, B2 => 
                           n22857, ZN => n3841);
   U14613 : OAI22_X1 port map( A1 => n16637, A2 => n23583, B1 => n20256, B2 => 
                           n22857, ZN => n3842);
   U14614 : OAI22_X1 port map( A1 => n16660, A2 => n23534, B1 => n20599, B2 => 
                           n22825, ZN => n3499);
   U14615 : OAI22_X1 port map( A1 => n16659, A2 => n23534, B1 => n20598, B2 => 
                           n22825, ZN => n3500);
   U14616 : OAI22_X1 port map( A1 => n16651, A2 => n23534, B1 => n20590, B2 => 
                           n22826, ZN => n3508);
   U14617 : OAI22_X1 port map( A1 => n16650, A2 => n23534, B1 => n20589, B2 => 
                           n22826, ZN => n3509);
   U14618 : OAI22_X1 port map( A1 => n16649, A2 => n23534, B1 => n20588, B2 => 
                           n22826, ZN => n3510);
   U14619 : OAI22_X1 port map( A1 => n16648, A2 => n23533, B1 => n20587, B2 => 
                           n22826, ZN => n3511);
   U14620 : OAI22_X1 port map( A1 => n16647, A2 => n23533, B1 => n20586, B2 => 
                           n22826, ZN => n3512);
   U14621 : OAI22_X1 port map( A1 => n16639, A2 => n23533, B1 => n20578, B2 => 
                           n22827, ZN => n3520);
   U14622 : OAI22_X1 port map( A1 => n16638, A2 => n23533, B1 => n20577, B2 => 
                           n22827, ZN => n3521);
   U14623 : OAI22_X1 port map( A1 => n16637, A2 => n23533, B1 => n20576, B2 => 
                           n22827, ZN => n3522);
   U14624 : OAI22_X1 port map( A1 => n16660, A2 => n23554, B1 => n20471, B2 => 
                           n22837, ZN => n3627);
   U14625 : OAI22_X1 port map( A1 => n16659, A2 => n23554, B1 => n20470, B2 => 
                           n22837, ZN => n3628);
   U14626 : OAI22_X1 port map( A1 => n16651, A2 => n23554, B1 => n20462, B2 => 
                           n22838, ZN => n3636);
   U14627 : OAI22_X1 port map( A1 => n16650, A2 => n23554, B1 => n20461, B2 => 
                           n22838, ZN => n3637);
   U14628 : OAI22_X1 port map( A1 => n16649, A2 => n23554, B1 => n20460, B2 => 
                           n22838, ZN => n3638);
   U14629 : OAI22_X1 port map( A1 => n16648, A2 => n23553, B1 => n20459, B2 => 
                           n22838, ZN => n3639);
   U14630 : OAI22_X1 port map( A1 => n16647, A2 => n23553, B1 => n20458, B2 => 
                           n22838, ZN => n3640);
   U14631 : OAI22_X1 port map( A1 => n16639, A2 => n23553, B1 => n20450, B2 => 
                           n22839, ZN => n3648);
   U14632 : OAI22_X1 port map( A1 => n16638, A2 => n23553, B1 => n20449, B2 => 
                           n22839, ZN => n3649);
   U14633 : OAI22_X1 port map( A1 => n16637, A2 => n23553, B1 => n20448, B2 => 
                           n22839, ZN => n3650);
   U14634 : OAI22_X1 port map( A1 => n16660, A2 => n23544, B1 => n20535, B2 => 
                           n22831, ZN => n3563);
   U14635 : OAI22_X1 port map( A1 => n16659, A2 => n23544, B1 => n20534, B2 => 
                           n22831, ZN => n3564);
   U14636 : OAI22_X1 port map( A1 => n16651, A2 => n23544, B1 => n20526, B2 => 
                           n22832, ZN => n3572);
   U14637 : OAI22_X1 port map( A1 => n16650, A2 => n23544, B1 => n20525, B2 => 
                           n22832, ZN => n3573);
   U14638 : OAI22_X1 port map( A1 => n16649, A2 => n23544, B1 => n20524, B2 => 
                           n22832, ZN => n3574);
   U14639 : OAI22_X1 port map( A1 => n16648, A2 => n23543, B1 => n20523, B2 => 
                           n22832, ZN => n3575);
   U14640 : OAI22_X1 port map( A1 => n16647, A2 => n23543, B1 => n20522, B2 => 
                           n22832, ZN => n3576);
   U14641 : OAI22_X1 port map( A1 => n16639, A2 => n23543, B1 => n20514, B2 => 
                           n22833, ZN => n3584);
   U14642 : OAI22_X1 port map( A1 => n16638, A2 => n23543, B1 => n20513, B2 => 
                           n22833, ZN => n3585);
   U14643 : OAI22_X1 port map( A1 => n16637, A2 => n23543, B1 => n20512, B2 => 
                           n22833, ZN => n3586);
   U14644 : OAI22_X1 port map( A1 => n16660, A2 => n23524, B1 => n20663, B2 => 
                           n22819, ZN => n3435);
   U14645 : OAI22_X1 port map( A1 => n16659, A2 => n23524, B1 => n20662, B2 => 
                           n22819, ZN => n3436);
   U14646 : OAI22_X1 port map( A1 => n16651, A2 => n23524, B1 => n20654, B2 => 
                           n22820, ZN => n3444);
   U14647 : OAI22_X1 port map( A1 => n16650, A2 => n23524, B1 => n20653, B2 => 
                           n22820, ZN => n3445);
   U14648 : OAI22_X1 port map( A1 => n16649, A2 => n23524, B1 => n20652, B2 => 
                           n22820, ZN => n3446);
   U14649 : OAI22_X1 port map( A1 => n16648, A2 => n23523, B1 => n20651, B2 => 
                           n22820, ZN => n3447);
   U14650 : OAI22_X1 port map( A1 => n16647, A2 => n23523, B1 => n20650, B2 => 
                           n22820, ZN => n3448);
   U14651 : OAI22_X1 port map( A1 => n16639, A2 => n23523, B1 => n20642, B2 => 
                           n22821, ZN => n3456);
   U14652 : OAI22_X1 port map( A1 => n16638, A2 => n23523, B1 => n20641, B2 => 
                           n22821, ZN => n3457);
   U14653 : OAI22_X1 port map( A1 => n16637, A2 => n23523, B1 => n20640, B2 => 
                           n22821, ZN => n3458);
   U14654 : OAI22_X1 port map( A1 => n16660, A2 => n23564, B1 => n20407, B2 => 
                           n22843, ZN => n3691);
   U14655 : OAI22_X1 port map( A1 => n16659, A2 => n23564, B1 => n20406, B2 => 
                           n22843, ZN => n3692);
   U14656 : OAI22_X1 port map( A1 => n16651, A2 => n23564, B1 => n20398, B2 => 
                           n22844, ZN => n3700);
   U14657 : OAI22_X1 port map( A1 => n16650, A2 => n23564, B1 => n20397, B2 => 
                           n22844, ZN => n3701);
   U14658 : OAI22_X1 port map( A1 => n16649, A2 => n23564, B1 => n20396, B2 => 
                           n22844, ZN => n3702);
   U14659 : OAI22_X1 port map( A1 => n16648, A2 => n23563, B1 => n20395, B2 => 
                           n22844, ZN => n3703);
   U14660 : OAI22_X1 port map( A1 => n16647, A2 => n23563, B1 => n20394, B2 => 
                           n22844, ZN => n3704);
   U14661 : OAI22_X1 port map( A1 => n16639, A2 => n23563, B1 => n20386, B2 => 
                           n22845, ZN => n3712);
   U14662 : OAI22_X1 port map( A1 => n16638, A2 => n23563, B1 => n20385, B2 => 
                           n22845, ZN => n3713);
   U14663 : OAI22_X1 port map( A1 => n16637, A2 => n23563, B1 => n20384, B2 => 
                           n22845, ZN => n3714);
   U14664 : OAI22_X1 port map( A1 => n16660, A2 => n23574, B1 => n20343, B2 => 
                           n22849, ZN => n3755);
   U14665 : OAI22_X1 port map( A1 => n16659, A2 => n23574, B1 => n20342, B2 => 
                           n22849, ZN => n3756);
   U14666 : OAI22_X1 port map( A1 => n16651, A2 => n23574, B1 => n20334, B2 => 
                           n22850, ZN => n3764);
   U14667 : OAI22_X1 port map( A1 => n16650, A2 => n23574, B1 => n20333, B2 => 
                           n22850, ZN => n3765);
   U14668 : OAI22_X1 port map( A1 => n16649, A2 => n23574, B1 => n20332, B2 => 
                           n22850, ZN => n3766);
   U14669 : OAI22_X1 port map( A1 => n16648, A2 => n23573, B1 => n20331, B2 => 
                           n22850, ZN => n3767);
   U14670 : OAI22_X1 port map( A1 => n16647, A2 => n23573, B1 => n20330, B2 => 
                           n22850, ZN => n3768);
   U14671 : OAI22_X1 port map( A1 => n16639, A2 => n23573, B1 => n20322, B2 => 
                           n22851, ZN => n3776);
   U14672 : OAI22_X1 port map( A1 => n16638, A2 => n23573, B1 => n20321, B2 => 
                           n22851, ZN => n3777);
   U14673 : OAI22_X1 port map( A1 => n16637, A2 => n23573, B1 => n20320, B2 => 
                           n22851, ZN => n3778);
   U14674 : OAI22_X1 port map( A1 => n16636, A2 => n23632, B1 => n19935, B2 => 
                           n22887, ZN => n4163);
   U14675 : OAI22_X1 port map( A1 => n16628, A2 => n23632, B1 => n19927, B2 => 
                           n22890, ZN => n4171);
   U14676 : OAI22_X1 port map( A1 => n16627, A2 => n23632, B1 => n19926, B2 => 
                           n22888, ZN => n4172);
   U14677 : OAI22_X1 port map( A1 => n16626, A2 => n23632, B1 => n19925, B2 => 
                           n22888, ZN => n4173);
   U14678 : OAI22_X1 port map( A1 => n16625, A2 => n23632, B1 => n19924, B2 => 
                           n22888, ZN => n4174);
   U14679 : OAI22_X1 port map( A1 => n16624, A2 => n23633, B1 => n19923, B2 => 
                           n22888, ZN => n4175);
   U14680 : OAI22_X1 port map( A1 => n16616, A2 => n23632, B1 => n19915, B2 => 
                           n22888, ZN => n4183);
   U14681 : OAI22_X1 port map( A1 => n16615, A2 => n23634, B1 => n19914, B2 => 
                           n22889, ZN => n4184);
   U14682 : OAI22_X1 port map( A1 => n16614, A2 => n23633, B1 => n19913, B2 => 
                           n22889, ZN => n4185);
   U14683 : OAI22_X1 port map( A1 => n16613, A2 => n23632, B1 => n19912, B2 => 
                           n22889, ZN => n4186);
   U14684 : OAI22_X1 port map( A1 => n16612, A2 => n23633, B1 => n19911, B2 => 
                           n22889, ZN => n4187);
   U14685 : OAI22_X1 port map( A1 => n16604, A2 => n23632, B1 => n19903, B2 => 
                           n22889, ZN => n4195);
   U14686 : OAI22_X1 port map( A1 => n16603, A2 => n23634, B1 => n19902, B2 => 
                           n22890, ZN => n4196);
   U14687 : OAI22_X1 port map( A1 => n16602, A2 => n23634, B1 => n19901, B2 => 
                           n22890, ZN => n4197);
   U14688 : OAI22_X1 port map( A1 => n16601, A2 => n23633, B1 => n19900, B2 => 
                           n22890, ZN => n4198);
   U14689 : OAI22_X1 port map( A1 => n16636, A2 => n23592, B1 => n20191, B2 => 
                           n22863, ZN => n3907);
   U14690 : OAI22_X1 port map( A1 => n16628, A2 => n23592, B1 => n20183, B2 => 
                           n22866, ZN => n3915);
   U14691 : OAI22_X1 port map( A1 => n16627, A2 => n23592, B1 => n20182, B2 => 
                           n22864, ZN => n3916);
   U14692 : OAI22_X1 port map( A1 => n16626, A2 => n23592, B1 => n20181, B2 => 
                           n22864, ZN => n3917);
   U14693 : OAI22_X1 port map( A1 => n16625, A2 => n23592, B1 => n20180, B2 => 
                           n22864, ZN => n3918);
   U14694 : OAI22_X1 port map( A1 => n16624, A2 => n23593, B1 => n20179, B2 => 
                           n22864, ZN => n3919);
   U14695 : OAI22_X1 port map( A1 => n16616, A2 => n23592, B1 => n20171, B2 => 
                           n22864, ZN => n3927);
   U14696 : OAI22_X1 port map( A1 => n16615, A2 => n23594, B1 => n20170, B2 => 
                           n22865, ZN => n3928);
   U14697 : OAI22_X1 port map( A1 => n16614, A2 => n23593, B1 => n20169, B2 => 
                           n22865, ZN => n3929);
   U14698 : OAI22_X1 port map( A1 => n16613, A2 => n23592, B1 => n20168, B2 => 
                           n22865, ZN => n3930);
   U14699 : OAI22_X1 port map( A1 => n16612, A2 => n23593, B1 => n20167, B2 => 
                           n22865, ZN => n3931);
   U14700 : OAI22_X1 port map( A1 => n16604, A2 => n23592, B1 => n20159, B2 => 
                           n22865, ZN => n3939);
   U14701 : OAI22_X1 port map( A1 => n16603, A2 => n23594, B1 => n20158, B2 => 
                           n22866, ZN => n3940);
   U14702 : OAI22_X1 port map( A1 => n16602, A2 => n23594, B1 => n20157, B2 => 
                           n22866, ZN => n3941);
   U14703 : OAI22_X1 port map( A1 => n16601, A2 => n23593, B1 => n20156, B2 => 
                           n22866, ZN => n3942);
   U14704 : OAI22_X1 port map( A1 => n16636, A2 => n23612, B1 => n20063, B2 => 
                           n22875, ZN => n4035);
   U14705 : OAI22_X1 port map( A1 => n16628, A2 => n23612, B1 => n20055, B2 => 
                           n22878, ZN => n4043);
   U14706 : OAI22_X1 port map( A1 => n16627, A2 => n23612, B1 => n20054, B2 => 
                           n22876, ZN => n4044);
   U14707 : OAI22_X1 port map( A1 => n16626, A2 => n23612, B1 => n20053, B2 => 
                           n22876, ZN => n4045);
   U14708 : OAI22_X1 port map( A1 => n16625, A2 => n23612, B1 => n20052, B2 => 
                           n22876, ZN => n4046);
   U14709 : OAI22_X1 port map( A1 => n16624, A2 => n23613, B1 => n20051, B2 => 
                           n22876, ZN => n4047);
   U14710 : OAI22_X1 port map( A1 => n16616, A2 => n23612, B1 => n20043, B2 => 
                           n22876, ZN => n4055);
   U14711 : OAI22_X1 port map( A1 => n16615, A2 => n23614, B1 => n20042, B2 => 
                           n22877, ZN => n4056);
   U14712 : OAI22_X1 port map( A1 => n16614, A2 => n23613, B1 => n20041, B2 => 
                           n22877, ZN => n4057);
   U14713 : OAI22_X1 port map( A1 => n16613, A2 => n23612, B1 => n20040, B2 => 
                           n22877, ZN => n4058);
   U14714 : OAI22_X1 port map( A1 => n16612, A2 => n23613, B1 => n20039, B2 => 
                           n22877, ZN => n4059);
   U14715 : OAI22_X1 port map( A1 => n16604, A2 => n23612, B1 => n20031, B2 => 
                           n22877, ZN => n4067);
   U14716 : OAI22_X1 port map( A1 => n16603, A2 => n23614, B1 => n20030, B2 => 
                           n22878, ZN => n4068);
   U14717 : OAI22_X1 port map( A1 => n16602, A2 => n23614, B1 => n20029, B2 => 
                           n22878, ZN => n4069);
   U14718 : OAI22_X1 port map( A1 => n16601, A2 => n23613, B1 => n20028, B2 => 
                           n22878, ZN => n4070);
   U14719 : OAI22_X1 port map( A1 => n16664, A2 => n23584, B1 => n20283, B2 => 
                           n22855, ZN => n3815);
   U14720 : OAI22_X1 port map( A1 => n16663, A2 => n23583, B1 => n20282, B2 => 
                           n22855, ZN => n3816);
   U14721 : OAI22_X1 port map( A1 => n16662, A2 => n23584, B1 => n20281, B2 => 
                           n22855, ZN => n3817);
   U14722 : OAI22_X1 port map( A1 => n16661, A2 => n23583, B1 => n20280, B2 => 
                           n22855, ZN => n3818);
   U14723 : OAI22_X1 port map( A1 => n16664, A2 => n23534, B1 => n20603, B2 => 
                           n22825, ZN => n3495);
   U14724 : OAI22_X1 port map( A1 => n16663, A2 => n23533, B1 => n20602, B2 => 
                           n22825, ZN => n3496);
   U14725 : OAI22_X1 port map( A1 => n16662, A2 => n23534, B1 => n20601, B2 => 
                           n22825, ZN => n3497);
   U14726 : OAI22_X1 port map( A1 => n16661, A2 => n23533, B1 => n20600, B2 => 
                           n22825, ZN => n3498);
   U14727 : OAI22_X1 port map( A1 => n16664, A2 => n23554, B1 => n20475, B2 => 
                           n22837, ZN => n3623);
   U14728 : OAI22_X1 port map( A1 => n16663, A2 => n23553, B1 => n20474, B2 => 
                           n22837, ZN => n3624);
   U14729 : OAI22_X1 port map( A1 => n16662, A2 => n23554, B1 => n20473, B2 => 
                           n22837, ZN => n3625);
   U14730 : OAI22_X1 port map( A1 => n16661, A2 => n23553, B1 => n20472, B2 => 
                           n22837, ZN => n3626);
   U14731 : OAI22_X1 port map( A1 => n16664, A2 => n23544, B1 => n20539, B2 => 
                           n22831, ZN => n3559);
   U14732 : OAI22_X1 port map( A1 => n16663, A2 => n23543, B1 => n20538, B2 => 
                           n22831, ZN => n3560);
   U14733 : OAI22_X1 port map( A1 => n16662, A2 => n23544, B1 => n20537, B2 => 
                           n22831, ZN => n3561);
   U14734 : OAI22_X1 port map( A1 => n16661, A2 => n23543, B1 => n20536, B2 => 
                           n22831, ZN => n3562);
   U14735 : OAI22_X1 port map( A1 => n16664, A2 => n23524, B1 => n20667, B2 => 
                           n22819, ZN => n3431);
   U14736 : OAI22_X1 port map( A1 => n16663, A2 => n23523, B1 => n20666, B2 => 
                           n22819, ZN => n3432);
   U14737 : OAI22_X1 port map( A1 => n16662, A2 => n23524, B1 => n20665, B2 => 
                           n22819, ZN => n3433);
   U14738 : OAI22_X1 port map( A1 => n16661, A2 => n23523, B1 => n20664, B2 => 
                           n22819, ZN => n3434);
   U14739 : OAI22_X1 port map( A1 => n16664, A2 => n23564, B1 => n20411, B2 => 
                           n22843, ZN => n3687);
   U14740 : OAI22_X1 port map( A1 => n16663, A2 => n23563, B1 => n20410, B2 => 
                           n22843, ZN => n3688);
   U14741 : OAI22_X1 port map( A1 => n16662, A2 => n23564, B1 => n20409, B2 => 
                           n22843, ZN => n3689);
   U14742 : OAI22_X1 port map( A1 => n16661, A2 => n23563, B1 => n20408, B2 => 
                           n22843, ZN => n3690);
   U14743 : OAI22_X1 port map( A1 => n16664, A2 => n23574, B1 => n20347, B2 => 
                           n22849, ZN => n3751);
   U14744 : OAI22_X1 port map( A1 => n16663, A2 => n23573, B1 => n20346, B2 => 
                           n22849, ZN => n3752);
   U14745 : OAI22_X1 port map( A1 => n16662, A2 => n23574, B1 => n20345, B2 => 
                           n22849, ZN => n3753);
   U14746 : OAI22_X1 port map( A1 => n16661, A2 => n23573, B1 => n20344, B2 => 
                           n22849, ZN => n3754);
   U14747 : AOI221_X1 port map( B1 => n23874, B2 => n21227, C1 => n23858, C2 =>
                           n21712, A => n15279, ZN => n15278);
   U14748 : OAI22_X1 port map( A1 => n18974, A2 => n23314, B1 => n19102, B2 => 
                           n23326, ZN => n15279);
   U14749 : AOI221_X1 port map( B1 => n23874, B2 => n21226, C1 => n23858, C2 =>
                           n21711, A => n15258, ZN => n15257);
   U14750 : OAI22_X1 port map( A1 => n18970, A2 => n23314, B1 => n19098, B2 => 
                           n23326, ZN => n15258);
   U14751 : AOI221_X1 port map( B1 => n23874, B2 => n21225, C1 => n23858, C2 =>
                           n21710, A => n15237, ZN => n15236);
   U14752 : OAI22_X1 port map( A1 => n18973, A2 => n23310, B1 => n19101, B2 => 
                           n23326, ZN => n15237);
   U14753 : AOI221_X1 port map( B1 => n23865, B2 => n21210, C1 => n23849, C2 =>
                           n21695, A => n15197, ZN => n15193);
   U14754 : OAI22_X1 port map( A1 => n18971, A2 => n23314, B1 => n19099, B2 => 
                           n23326, ZN => n15197);
   U14755 : AOI221_X1 port map( B1 => n23842, B2 => n21829, C1 => n23816, C2 =>
                           n22144, A => n15280, ZN => n15277);
   U14756 : OAI22_X1 port map( A1 => n18782, A2 => n23286, B1 => n18910, B2 => 
                           n23303, ZN => n15280);
   U14757 : AOI221_X1 port map( B1 => n23842, B2 => n21828, C1 => n23816, C2 =>
                           n22038, A => n15259, ZN => n15256);
   U14758 : OAI22_X1 port map( A1 => n18778, A2 => n23291, B1 => n18906, B2 => 
                           n23303, ZN => n15259);
   U14759 : AOI221_X1 port map( B1 => n23842, B2 => n21827, C1 => n23816, C2 =>
                           n22037, A => n15238, ZN => n15235);
   U14760 : OAI22_X1 port map( A1 => n18781, A2 => n23287, B1 => n18909, B2 => 
                           n23303, ZN => n15238);
   U14761 : AOI221_X1 port map( B1 => n23833, B2 => n21826, C1 => n23816, C2 =>
                           n22143, A => n15200, ZN => n15192);
   U14762 : OAI22_X1 port map( A1 => n18779, A2 => n23291, B1 => n18907, B2 => 
                           n23303, ZN => n15200);
   U14763 : AOI221_X1 port map( B1 => n23872, B2 => n21232, C1 => n23856, C2 =>
                           n21717, A => n15531, ZN => n15530);
   U14764 : OAI22_X1 port map( A1 => n18980, A2 => n23311, B1 => n19108, B2 => 
                           n23325, ZN => n15531);
   U14765 : AOI221_X1 port map( B1 => n23872, B2 => n21279, C1 => n23856, C2 =>
                           n21835, A => n15510, ZN => n15509);
   U14766 : OAI22_X1 port map( A1 => n18964, A2 => n23312, B1 => n19092, B2 => 
                           n23325, ZN => n15510);
   U14767 : AOI221_X1 port map( B1 => n23873, B2 => n21231, C1 => n23857, C2 =>
                           n21716, A => n15489, ZN => n15488);
   U14768 : OAI22_X1 port map( A1 => n18979, A2 => n23313, B1 => n19107, B2 => 
                           n23325, ZN => n15489);
   U14769 : AOI221_X1 port map( B1 => n23873, B2 => n21247, C1 => n23857, C2 =>
                           n21731, A => n15468, ZN => n15467);
   U14770 : OAI22_X1 port map( A1 => n18965, A2 => n23314, B1 => n19093, B2 => 
                           n23325, ZN => n15468);
   U14771 : AOI221_X1 port map( B1 => n23873, B2 => n21230, C1 => n23857, C2 =>
                           n21715, A => n15447, ZN => n15446);
   U14772 : OAI22_X1 port map( A1 => n18978, A2 => n23310, B1 => n19106, B2 => 
                           n23325, ZN => n15447);
   U14773 : AOI221_X1 port map( B1 => n23873, B2 => n21229, C1 => n23857, C2 =>
                           n21714, A => n15426, ZN => n15425);
   U14774 : OAI22_X1 port map( A1 => n18966, A2 => n23309, B1 => n19094, B2 => 
                           n23325, ZN => n15426);
   U14775 : AOI221_X1 port map( B1 => n23873, B2 => n21246, C1 => n23857, C2 =>
                           n21730, A => n15405, ZN => n15404);
   U14776 : OAI22_X1 port map( A1 => n18977, A2 => n23314, B1 => n19105, B2 => 
                           n23326, ZN => n15405);
   U14777 : AOI221_X1 port map( B1 => n23873, B2 => n21266, C1 => n23857, C2 =>
                           n21754, A => n15384, ZN => n15383);
   U14778 : OAI22_X1 port map( A1 => n18967, A2 => n23314, B1 => n19095, B2 => 
                           n23326, ZN => n15384);
   U14779 : AOI221_X1 port map( B1 => n23873, B2 => n21245, C1 => n23857, C2 =>
                           n21729, A => n15363, ZN => n15362);
   U14780 : OAI22_X1 port map( A1 => n18976, A2 => n23314, B1 => n19104, B2 => 
                           n23326, ZN => n15363);
   U14781 : AOI221_X1 port map( B1 => n23874, B2 => n21244, C1 => n23858, C2 =>
                           n21728, A => n15342, ZN => n15341);
   U14782 : OAI22_X1 port map( A1 => n18968, A2 => n23314, B1 => n19096, B2 => 
                           n23326, ZN => n15342);
   U14783 : AOI221_X1 port map( B1 => n23874, B2 => n21228, C1 => n23858, C2 =>
                           n21713, A => n15321, ZN => n15320);
   U14784 : OAI22_X1 port map( A1 => n18975, A2 => n23314, B1 => n19103, B2 => 
                           n23325, ZN => n15321);
   U14785 : AOI221_X1 port map( B1 => n23874, B2 => n21211, C1 => n23858, C2 =>
                           n21696, A => n15300, ZN => n15299);
   U14786 : OAI22_X1 port map( A1 => n18969, A2 => n23314, B1 => n19097, B2 => 
                           n23326, ZN => n15300);
   U14787 : AOI221_X1 port map( B1 => n23840, B2 => n21778, C1 => n23818, C2 =>
                           n22154, A => n15532, ZN => n15529);
   U14788 : OAI22_X1 port map( A1 => n18788, A2 => n23288, B1 => n18916, B2 => 
                           n23302, ZN => n15532);
   U14789 : AOI221_X1 port map( B1 => n23840, B2 => n21777, C1 => n23818, C2 =>
                           n22040, A => n15511, ZN => n15508);
   U14790 : OAI22_X1 port map( A1 => n18772, A2 => n23289, B1 => n18900, B2 => 
                           n23302, ZN => n15511);
   U14791 : AOI221_X1 port map( B1 => n23841, B2 => n21776, C1 => n23818, C2 =>
                           n22153, A => n15490, ZN => n15487);
   U14792 : OAI22_X1 port map( A1 => n18787, A2 => n23290, B1 => n18915, B2 => 
                           n23302, ZN => n15490);
   U14793 : AOI221_X1 port map( B1 => n23841, B2 => n21775, C1 => n23818, C2 =>
                           n22152, A => n15469, ZN => n15466);
   U14794 : OAI22_X1 port map( A1 => n18773, A2 => n23286, B1 => n18901, B2 => 
                           n23302, ZN => n15469);
   U14795 : AOI221_X1 port map( B1 => n23841, B2 => n21774, C1 => n23817, C2 =>
                           n22151, A => n15448, ZN => n15445);
   U14796 : OAI22_X1 port map( A1 => n18786, A2 => n23287, B1 => n18914, B2 => 
                           n23302, ZN => n15448);
   U14797 : AOI221_X1 port map( B1 => n23841, B2 => n21773, C1 => n23817, C2 =>
                           n22150, A => n15427, ZN => n15424);
   U14798 : OAI22_X1 port map( A1 => n18774, A2 => n23291, B1 => n18902, B2 => 
                           n23302, ZN => n15427);
   U14799 : AOI221_X1 port map( B1 => n23841, B2 => n21772, C1 => n23817, C2 =>
                           n22149, A => n15406, ZN => n15403);
   U14800 : OAI22_X1 port map( A1 => n18785, A2 => n23291, B1 => n18913, B2 => 
                           n23303, ZN => n15406);
   U14801 : AOI221_X1 port map( B1 => n23841, B2 => n21771, C1 => n23817, C2 =>
                           n22039, A => n15385, ZN => n15382);
   U14802 : OAI22_X1 port map( A1 => n18775, A2 => n23291, B1 => n18903, B2 => 
                           n23303, ZN => n15385);
   U14803 : AOI221_X1 port map( B1 => n23841, B2 => n21770, C1 => n23817, C2 =>
                           n22148, A => n15364, ZN => n15361);
   U14804 : OAI22_X1 port map( A1 => n18784, A2 => n23291, B1 => n18912, B2 => 
                           n23303, ZN => n15364);
   U14805 : AOI221_X1 port map( B1 => n23842, B2 => n21769, C1 => n23817, C2 =>
                           n22147, A => n15343, ZN => n15340);
   U14806 : OAI22_X1 port map( A1 => n18776, A2 => n23291, B1 => n18904, B2 => 
                           n23303, ZN => n15343);
   U14807 : AOI221_X1 port map( B1 => n23842, B2 => n21768, C1 => n23816, C2 =>
                           n22146, A => n15322, ZN => n15319);
   U14808 : OAI22_X1 port map( A1 => n18783, A2 => n23291, B1 => n18911, B2 => 
                           n23302, ZN => n15322);
   U14809 : AOI221_X1 port map( B1 => n23842, B2 => n21767, C1 => n23816, C2 =>
                           n22145, A => n15301, ZN => n15298);
   U14810 : OAI22_X1 port map( A1 => n18777, A2 => n23291, B1 => n18905, B2 => 
                           n23303, ZN => n15301);
   U14811 : AOI221_X1 port map( B1 => n23842, B2 => n22379, C1 => n23816, C2 =>
                           n22304, A => n15284, ZN => n15281);
   U14812 : OAI22_X1 port map( A1 => n19294, A2 => n23291, B1 => n19422, B2 => 
                           n23303, ZN => n15284);
   U14813 : AOI221_X1 port map( B1 => n23842, B2 => n22324, C1 => n23816, C2 =>
                           n22345, A => n15263, ZN => n15260);
   U14814 : OAI22_X1 port map( A1 => n19290, A2 => n23291, B1 => n19418, B2 => 
                           n23303, ZN => n15263);
   U14815 : AOI221_X1 port map( B1 => n23842, B2 => n22326, C1 => n23816, C2 =>
                           n22303, A => n15242, ZN => n15239);
   U14816 : OAI22_X1 port map( A1 => n19293, A2 => n23288, B1 => n19421, B2 => 
                           n23303, ZN => n15242);
   U14817 : AOI221_X1 port map( B1 => n23842, B2 => n22325, C1 => n23816, C2 =>
                           n22302, A => n15205, ZN => n15201);
   U14818 : OAI22_X1 port map( A1 => n19291, A2 => n23291, B1 => n19419, B2 => 
                           n23303, ZN => n15205);
   U14819 : AOI221_X1 port map( B1 => n23874, B2 => n21183, C1 => n23858, C2 =>
                           n21596, A => n15283, ZN => n15282);
   U14820 : OAI22_X1 port map( A1 => n19486, A2 => n23309, B1 => n19614, B2 => 
                           n23326, ZN => n15283);
   U14821 : AOI221_X1 port map( B1 => n23874, B2 => n21158, C1 => n23858, C2 =>
                           n21595, A => n15262, ZN => n15261);
   U14822 : OAI22_X1 port map( A1 => n19482, A2 => n23314, B1 => n19610, B2 => 
                           n23326, ZN => n15262);
   U14823 : AOI221_X1 port map( B1 => n23874, B2 => n21182, C1 => n23858, C2 =>
                           n21594, A => n15241, ZN => n15240);
   U14824 : OAI22_X1 port map( A1 => n19485, A2 => n23311, B1 => n19613, B2 => 
                           n23326, ZN => n15241);
   U14825 : AOI221_X1 port map( B1 => n23874, B2 => n21151, C1 => n23858, C2 =>
                           n21579, A => n15204, ZN => n15202);
   U14826 : OAI22_X1 port map( A1 => n19483, A2 => n23314, B1 => n19611, B2 => 
                           n23326, ZN => n15204);
   U14827 : OAI22_X1 port map( A1 => n16658, A2 => n23604, B1 => n20149, B2 => 
                           n22867, ZN => n3949);
   U14828 : OAI22_X1 port map( A1 => n16657, A2 => n23604, B1 => n20148, B2 => 
                           n22867, ZN => n3950);
   U14829 : OAI22_X1 port map( A1 => n16656, A2 => n23604, B1 => n20147, B2 => 
                           n22867, ZN => n3951);
   U14830 : OAI22_X1 port map( A1 => n16655, A2 => n23604, B1 => n20146, B2 => 
                           n22867, ZN => n3952);
   U14831 : OAI22_X1 port map( A1 => n16654, A2 => n23604, B1 => n20145, B2 => 
                           n22867, ZN => n3953);
   U14832 : OAI22_X1 port map( A1 => n16653, A2 => n23604, B1 => n20144, B2 => 
                           n22867, ZN => n3954);
   U14833 : OAI22_X1 port map( A1 => n16652, A2 => n23604, B1 => n20143, B2 => 
                           n22868, ZN => n3955);
   U14834 : OAI22_X1 port map( A1 => n16646, A2 => n23603, B1 => n20137, B2 => 
                           n22868, ZN => n3961);
   U14835 : OAI22_X1 port map( A1 => n16645, A2 => n23603, B1 => n20136, B2 => 
                           n22868, ZN => n3962);
   U14836 : OAI22_X1 port map( A1 => n16644, A2 => n23603, B1 => n20135, B2 => 
                           n22868, ZN => n3963);
   U14837 : OAI22_X1 port map( A1 => n16643, A2 => n23603, B1 => n20134, B2 => 
                           n22868, ZN => n3964);
   U14838 : OAI22_X1 port map( A1 => n16642, A2 => n23603, B1 => n20133, B2 => 
                           n22868, ZN => n3965);
   U14839 : OAI22_X1 port map( A1 => n16641, A2 => n23603, B1 => n20132, B2 => 
                           n22868, ZN => n3966);
   U14840 : OAI22_X1 port map( A1 => n16640, A2 => n23603, B1 => n20131, B2 => 
                           n22869, ZN => n3967);
   U14841 : OAI22_X1 port map( A1 => n16658, A2 => n23624, B1 => n20021, B2 => 
                           n22879, ZN => n4077);
   U14842 : OAI22_X1 port map( A1 => n16657, A2 => n23624, B1 => n20020, B2 => 
                           n22879, ZN => n4078);
   U14843 : OAI22_X1 port map( A1 => n16656, A2 => n23624, B1 => n20019, B2 => 
                           n22879, ZN => n4079);
   U14844 : OAI22_X1 port map( A1 => n16655, A2 => n23624, B1 => n20018, B2 => 
                           n22879, ZN => n4080);
   U14845 : OAI22_X1 port map( A1 => n16654, A2 => n23624, B1 => n20017, B2 => 
                           n22879, ZN => n4081);
   U14846 : OAI22_X1 port map( A1 => n16653, A2 => n23624, B1 => n20016, B2 => 
                           n22879, ZN => n4082);
   U14847 : OAI22_X1 port map( A1 => n16652, A2 => n23624, B1 => n20015, B2 => 
                           n22880, ZN => n4083);
   U14848 : OAI22_X1 port map( A1 => n16646, A2 => n23623, B1 => n20009, B2 => 
                           n22880, ZN => n4089);
   U14849 : OAI22_X1 port map( A1 => n16645, A2 => n23623, B1 => n20008, B2 => 
                           n22880, ZN => n4090);
   U14850 : OAI22_X1 port map( A1 => n16644, A2 => n23623, B1 => n20007, B2 => 
                           n22880, ZN => n4091);
   U14851 : OAI22_X1 port map( A1 => n16643, A2 => n23623, B1 => n20006, B2 => 
                           n22880, ZN => n4092);
   U14852 : OAI22_X1 port map( A1 => n16642, A2 => n23623, B1 => n20005, B2 => 
                           n22880, ZN => n4093);
   U14853 : OAI22_X1 port map( A1 => n16641, A2 => n23623, B1 => n20004, B2 => 
                           n22880, ZN => n4094);
   U14854 : OAI22_X1 port map( A1 => n16640, A2 => n23623, B1 => n20003, B2 => 
                           n22881, ZN => n4095);
   U14855 : OAI22_X1 port map( A1 => n16658, A2 => n23644, B1 => n19893, B2 => 
                           n22891, ZN => n4205);
   U14856 : OAI22_X1 port map( A1 => n16657, A2 => n23644, B1 => n19892, B2 => 
                           n22891, ZN => n4206);
   U14857 : OAI22_X1 port map( A1 => n16656, A2 => n23644, B1 => n19891, B2 => 
                           n22891, ZN => n4207);
   U14858 : OAI22_X1 port map( A1 => n16655, A2 => n23644, B1 => n19890, B2 => 
                           n22891, ZN => n4208);
   U14859 : OAI22_X1 port map( A1 => n16654, A2 => n23644, B1 => n19889, B2 => 
                           n22891, ZN => n4209);
   U14860 : OAI22_X1 port map( A1 => n16653, A2 => n23644, B1 => n19888, B2 => 
                           n22891, ZN => n4210);
   U14861 : OAI22_X1 port map( A1 => n16652, A2 => n23644, B1 => n19887, B2 => 
                           n22892, ZN => n4211);
   U14862 : OAI22_X1 port map( A1 => n16646, A2 => n23643, B1 => n19881, B2 => 
                           n22892, ZN => n4217);
   U14863 : OAI22_X1 port map( A1 => n16645, A2 => n23643, B1 => n19880, B2 => 
                           n22892, ZN => n4218);
   U14864 : OAI22_X1 port map( A1 => n16644, A2 => n23643, B1 => n19879, B2 => 
                           n22892, ZN => n4219);
   U14865 : OAI22_X1 port map( A1 => n16643, A2 => n23643, B1 => n19878, B2 => 
                           n22892, ZN => n4220);
   U14866 : OAI22_X1 port map( A1 => n16642, A2 => n23643, B1 => n19877, B2 => 
                           n22892, ZN => n4221);
   U14867 : OAI22_X1 port map( A1 => n16641, A2 => n23643, B1 => n19876, B2 => 
                           n22892, ZN => n4222);
   U14868 : OAI22_X1 port map( A1 => n16640, A2 => n23643, B1 => n19875, B2 => 
                           n22893, ZN => n4223);
   U14869 : OAI22_X1 port map( A1 => n16658, A2 => n23664, B1 => n19765, B2 => 
                           n22903, ZN => n4333);
   U14870 : OAI22_X1 port map( A1 => n16657, A2 => n23664, B1 => n19764, B2 => 
                           n22903, ZN => n4334);
   U14871 : OAI22_X1 port map( A1 => n16656, A2 => n23664, B1 => n19763, B2 => 
                           n22903, ZN => n4335);
   U14872 : OAI22_X1 port map( A1 => n16655, A2 => n23664, B1 => n19762, B2 => 
                           n22903, ZN => n4336);
   U14873 : OAI22_X1 port map( A1 => n16654, A2 => n23664, B1 => n19761, B2 => 
                           n22903, ZN => n4337);
   U14874 : OAI22_X1 port map( A1 => n16653, A2 => n23664, B1 => n19760, B2 => 
                           n22903, ZN => n4338);
   U14875 : OAI22_X1 port map( A1 => n16652, A2 => n23664, B1 => n19759, B2 => 
                           n22904, ZN => n4339);
   U14876 : OAI22_X1 port map( A1 => n16646, A2 => n23663, B1 => n19753, B2 => 
                           n22904, ZN => n4345);
   U14877 : OAI22_X1 port map( A1 => n16645, A2 => n23663, B1 => n19752, B2 => 
                           n22904, ZN => n4346);
   U14878 : OAI22_X1 port map( A1 => n16644, A2 => n23663, B1 => n19751, B2 => 
                           n22904, ZN => n4347);
   U14879 : OAI22_X1 port map( A1 => n16643, A2 => n23663, B1 => n19750, B2 => 
                           n22904, ZN => n4348);
   U14880 : OAI22_X1 port map( A1 => n16642, A2 => n23663, B1 => n19749, B2 => 
                           n22904, ZN => n4349);
   U14881 : OAI22_X1 port map( A1 => n16641, A2 => n23663, B1 => n19748, B2 => 
                           n22904, ZN => n4350);
   U14882 : OAI22_X1 port map( A1 => n16640, A2 => n23663, B1 => n19747, B2 => 
                           n22905, ZN => n4351);
   U14883 : AOI221_X1 port map( B1 => n23840, B2 => n22327, C1 => n23818, C2 =>
                           n22357, A => n15536, ZN => n15533);
   U14884 : OAI22_X1 port map( A1 => n19300, A2 => n23290, B1 => n19428, B2 => 
                           n23302, ZN => n15536);
   U14885 : AOI221_X1 port map( B1 => n23840, B2 => n22388, C1 => n23818, C2 =>
                           n22348, A => n15515, ZN => n15512);
   U14886 : OAI22_X1 port map( A1 => n19284, A2 => n23286, B1 => n19412, B2 => 
                           n23302, ZN => n15515);
   U14887 : AOI221_X1 port map( B1 => n23840, B2 => n22395, C1 => n23818, C2 =>
                           n22356, A => n15494, ZN => n15491);
   U14888 : OAI22_X1 port map( A1 => n19299, A2 => n23287, B1 => n19427, B2 => 
                           n23302, ZN => n15494);
   U14889 : AOI221_X1 port map( B1 => n23840, B2 => n22402, C1 => n23818, C2 =>
                           n22349, A => n15473, ZN => n15470);
   U14890 : OAI22_X1 port map( A1 => n19285, A2 => n23291, B1 => n19413, B2 => 
                           n23302, ZN => n15473);
   U14891 : AOI221_X1 port map( B1 => n23841, B2 => n22394, C1 => n23817, C2 =>
                           n22355, A => n15452, ZN => n15449);
   U14892 : OAI22_X1 port map( A1 => n19298, A2 => n23288, B1 => n19426, B2 => 
                           n23302, ZN => n15452);
   U14893 : AOI221_X1 port map( B1 => n23841, B2 => n22389, C1 => n23817, C2 =>
                           n22350, A => n15431, ZN => n15428);
   U14894 : OAI22_X1 port map( A1 => n19286, A2 => n23289, B1 => n19414, B2 => 
                           n23302, ZN => n15431);
   U14895 : AOI221_X1 port map( B1 => n23841, B2 => n22393, C1 => n23817, C2 =>
                           n22360, A => n15410, ZN => n15407);
   U14896 : OAI22_X1 port map( A1 => n19297, A2 => n23291, B1 => n19425, B2 => 
                           n23302, ZN => n15410);
   U14897 : AOI221_X1 port map( B1 => n23841, B2 => n22390, C1 => n23817, C2 =>
                           n22351, A => n15389, ZN => n15386);
   U14898 : OAI22_X1 port map( A1 => n19287, A2 => n23291, B1 => n19415, B2 => 
                           n23303, ZN => n15389);
   U14899 : AOI221_X1 port map( B1 => n23841, B2 => n22392, C1 => n23817, C2 =>
                           n22354, A => n15368, ZN => n15365);
   U14900 : OAI22_X1 port map( A1 => n19296, A2 => n23291, B1 => n19424, B2 => 
                           n23303, ZN => n15368);
   U14901 : AOI221_X1 port map( B1 => n23841, B2 => n22322, C1 => n23817, C2 =>
                           n22301, A => n15347, ZN => n15344);
   U14902 : OAI22_X1 port map( A1 => n19288, A2 => n23291, B1 => n19416, B2 => 
                           n23300, ZN => n15347);
   U14903 : AOI221_X1 port map( B1 => n23842, B2 => n22391, C1 => n23816, C2 =>
                           n22353, A => n15326, ZN => n15323);
   U14904 : OAI22_X1 port map( A1 => n19295, A2 => n23291, B1 => n19423, B2 => 
                           n23301, ZN => n15326);
   U14905 : AOI221_X1 port map( B1 => n23842, B2 => n22323, C1 => n23816, C2 =>
                           n22352, A => n15305, ZN => n15302);
   U14906 : OAI22_X1 port map( A1 => n19289, A2 => n23291, B1 => n19417, B2 => 
                           n23301, ZN => n15305);
   U14907 : AOI221_X1 port map( B1 => n23872, B2 => n21187, C1 => n23856, C2 =>
                           n21601, A => n15535, ZN => n15534);
   U14908 : OAI22_X1 port map( A1 => n19492, A2 => n23313, B1 => n19620, B2 => 
                           n23325, ZN => n15535);
   U14909 : AOI221_X1 port map( B1 => n23872, B2 => n21278, C1 => n23856, C2 =>
                           n21758, A => n15514, ZN => n15513);
   U14910 : OAI22_X1 port map( A1 => n19476, A2 => n23314, B1 => n19604, B2 => 
                           n23325, ZN => n15514);
   U14911 : AOI221_X1 port map( B1 => n23872, B2 => n21186, C1 => n23856, C2 =>
                           n21600, A => n15493, ZN => n15492);
   U14912 : OAI22_X1 port map( A1 => n19491, A2 => n23310, B1 => n19619, B2 => 
                           n23325, ZN => n15493);
   U14913 : AOI221_X1 port map( B1 => n23872, B2 => n21194, C1 => n23856, C2 =>
                           n21614, A => n15472, ZN => n15471);
   U14914 : OAI22_X1 port map( A1 => n19477, A2 => n23309, B1 => n19605, B2 => 
                           n23325, ZN => n15472);
   U14915 : AOI221_X1 port map( B1 => n23873, B2 => n21185, C1 => n23857, C2 =>
                           n21599, A => n15451, ZN => n15450);
   U14916 : OAI22_X1 port map( A1 => n19490, A2 => n23311, B1 => n19618, B2 => 
                           n23325, ZN => n15451);
   U14917 : AOI221_X1 port map( B1 => n23873, B2 => n21159, C1 => n23857, C2 =>
                           n21598, A => n15430, ZN => n15429);
   U14918 : OAI22_X1 port map( A1 => n19478, A2 => n23312, B1 => n19606, B2 => 
                           n23325, ZN => n15430);
   U14919 : AOI221_X1 port map( B1 => n23873, B2 => n21165, C1 => n23857, C2 =>
                           n21613, A => n15409, ZN => n15408);
   U14920 : OAI22_X1 port map( A1 => n19489, A2 => n23314, B1 => n19617, B2 => 
                           n23325, ZN => n15409);
   U14921 : AOI221_X1 port map( B1 => n23873, B2 => n21207, C1 => n23857, C2 =>
                           n21636, A => n15388, ZN => n15387);
   U14922 : OAI22_X1 port map( A1 => n19479, A2 => n23314, B1 => n19607, B2 => 
                           n23326, ZN => n15388);
   U14923 : AOI221_X1 port map( B1 => n23873, B2 => n21193, C1 => n23857, C2 =>
                           n21612, A => n15367, ZN => n15366);
   U14924 : OAI22_X1 port map( A1 => n19488, A2 => n23314, B1 => n19616, B2 => 
                           n23326, ZN => n15367);
   U14925 : AOI221_X1 port map( B1 => n23873, B2 => n21164, C1 => n23857, C2 =>
                           n21611, A => n15346, ZN => n15345);
   U14926 : OAI22_X1 port map( A1 => n19480, A2 => n23314, B1 => n19608, B2 => 
                           n23323, ZN => n15346);
   U14927 : AOI221_X1 port map( B1 => n23874, B2 => n21184, C1 => n23858, C2 =>
                           n21597, A => n15325, ZN => n15324);
   U14928 : OAI22_X1 port map( A1 => n19487, A2 => n23314, B1 => n19615, B2 => 
                           n23324, ZN => n15325);
   U14929 : AOI221_X1 port map( B1 => n23874, B2 => n21174, C1 => n23858, C2 =>
                           n21580, A => n15304, ZN => n15303);
   U14930 : OAI22_X1 port map( A1 => n19481, A2 => n23314, B1 => n19609, B2 => 
                           n23324, ZN => n15304);
   U14931 : OAI22_X1 port map( A1 => n16660, A2 => n23644, B1 => n19895, B2 => 
                           n22891, ZN => n4203);
   U14932 : OAI22_X1 port map( A1 => n16659, A2 => n23644, B1 => n19894, B2 => 
                           n22891, ZN => n4204);
   U14933 : OAI22_X1 port map( A1 => n16651, A2 => n23644, B1 => n19886, B2 => 
                           n22892, ZN => n4212);
   U14934 : OAI22_X1 port map( A1 => n16650, A2 => n23644, B1 => n19885, B2 => 
                           n22892, ZN => n4213);
   U14935 : OAI22_X1 port map( A1 => n16649, A2 => n23644, B1 => n19884, B2 => 
                           n22892, ZN => n4214);
   U14936 : OAI22_X1 port map( A1 => n16648, A2 => n23643, B1 => n19883, B2 => 
                           n22892, ZN => n4215);
   U14937 : OAI22_X1 port map( A1 => n16647, A2 => n23643, B1 => n19882, B2 => 
                           n22892, ZN => n4216);
   U14938 : OAI22_X1 port map( A1 => n16639, A2 => n23643, B1 => n19874, B2 => 
                           n22893, ZN => n4224);
   U14939 : OAI22_X1 port map( A1 => n16638, A2 => n23643, B1 => n19873, B2 => 
                           n22893, ZN => n4225);
   U14940 : OAI22_X1 port map( A1 => n16637, A2 => n23643, B1 => n19872, B2 => 
                           n22893, ZN => n4226);
   U14941 : OAI22_X1 port map( A1 => n16660, A2 => n23664, B1 => n19767, B2 => 
                           n22903, ZN => n4331);
   U14942 : OAI22_X1 port map( A1 => n16659, A2 => n23664, B1 => n19766, B2 => 
                           n22903, ZN => n4332);
   U14943 : OAI22_X1 port map( A1 => n16651, A2 => n23664, B1 => n19758, B2 => 
                           n22904, ZN => n4340);
   U14944 : OAI22_X1 port map( A1 => n16650, A2 => n23664, B1 => n19757, B2 => 
                           n22904, ZN => n4341);
   U14945 : OAI22_X1 port map( A1 => n16649, A2 => n23664, B1 => n19756, B2 => 
                           n22904, ZN => n4342);
   U14946 : OAI22_X1 port map( A1 => n16648, A2 => n23663, B1 => n19755, B2 => 
                           n22904, ZN => n4343);
   U14947 : OAI22_X1 port map( A1 => n16647, A2 => n23663, B1 => n19754, B2 => 
                           n22904, ZN => n4344);
   U14948 : OAI22_X1 port map( A1 => n16639, A2 => n23663, B1 => n19746, B2 => 
                           n22905, ZN => n4352);
   U14949 : OAI22_X1 port map( A1 => n16638, A2 => n23663, B1 => n19745, B2 => 
                           n22905, ZN => n4353);
   U14950 : OAI22_X1 port map( A1 => n16637, A2 => n23663, B1 => n19744, B2 => 
                           n22905, ZN => n4354);
   U14951 : OAI22_X1 port map( A1 => n16660, A2 => n23604, B1 => n20151, B2 => 
                           n22867, ZN => n3947);
   U14952 : OAI22_X1 port map( A1 => n16659, A2 => n23604, B1 => n20150, B2 => 
                           n22867, ZN => n3948);
   U14953 : OAI22_X1 port map( A1 => n16651, A2 => n23604, B1 => n20142, B2 => 
                           n22868, ZN => n3956);
   U14954 : OAI22_X1 port map( A1 => n16650, A2 => n23604, B1 => n20141, B2 => 
                           n22868, ZN => n3957);
   U14955 : OAI22_X1 port map( A1 => n16649, A2 => n23604, B1 => n20140, B2 => 
                           n22868, ZN => n3958);
   U14956 : OAI22_X1 port map( A1 => n16648, A2 => n23603, B1 => n20139, B2 => 
                           n22868, ZN => n3959);
   U14957 : OAI22_X1 port map( A1 => n16647, A2 => n23603, B1 => n20138, B2 => 
                           n22868, ZN => n3960);
   U14958 : OAI22_X1 port map( A1 => n16639, A2 => n23603, B1 => n20130, B2 => 
                           n22869, ZN => n3968);
   U14959 : OAI22_X1 port map( A1 => n16638, A2 => n23603, B1 => n20129, B2 => 
                           n22869, ZN => n3969);
   U14960 : OAI22_X1 port map( A1 => n16637, A2 => n23603, B1 => n20128, B2 => 
                           n22869, ZN => n3970);
   U14961 : OAI22_X1 port map( A1 => n16660, A2 => n23624, B1 => n20023, B2 => 
                           n22879, ZN => n4075);
   U14962 : OAI22_X1 port map( A1 => n16659, A2 => n23624, B1 => n20022, B2 => 
                           n22879, ZN => n4076);
   U14963 : OAI22_X1 port map( A1 => n16651, A2 => n23624, B1 => n20014, B2 => 
                           n22880, ZN => n4084);
   U14964 : OAI22_X1 port map( A1 => n16650, A2 => n23624, B1 => n20013, B2 => 
                           n22880, ZN => n4085);
   U14965 : OAI22_X1 port map( A1 => n16649, A2 => n23624, B1 => n20012, B2 => 
                           n22880, ZN => n4086);
   U14966 : OAI22_X1 port map( A1 => n16648, A2 => n23623, B1 => n20011, B2 => 
                           n22880, ZN => n4087);
   U14967 : OAI22_X1 port map( A1 => n16647, A2 => n23623, B1 => n20010, B2 => 
                           n22880, ZN => n4088);
   U14968 : OAI22_X1 port map( A1 => n16639, A2 => n23623, B1 => n20002, B2 => 
                           n22881, ZN => n4096);
   U14969 : OAI22_X1 port map( A1 => n16638, A2 => n23623, B1 => n20001, B2 => 
                           n22881, ZN => n4097);
   U14970 : OAI22_X1 port map( A1 => n16637, A2 => n23623, B1 => n20000, B2 => 
                           n22881, ZN => n4098);
   U14971 : OAI22_X1 port map( A1 => n16658, A2 => n23654, B1 => n19829, B2 => 
                           n22897, ZN => n4269);
   U14972 : OAI22_X1 port map( A1 => n16657, A2 => n23654, B1 => n19828, B2 => 
                           n22897, ZN => n4270);
   U14973 : OAI22_X1 port map( A1 => n16656, A2 => n23654, B1 => n19827, B2 => 
                           n22897, ZN => n4271);
   U14974 : OAI22_X1 port map( A1 => n16655, A2 => n23654, B1 => n19826, B2 => 
                           n22897, ZN => n4272);
   U14975 : OAI22_X1 port map( A1 => n16654, A2 => n23654, B1 => n19825, B2 => 
                           n22897, ZN => n4273);
   U14976 : OAI22_X1 port map( A1 => n16653, A2 => n23654, B1 => n19824, B2 => 
                           n22897, ZN => n4274);
   U14977 : OAI22_X1 port map( A1 => n16652, A2 => n23654, B1 => n19823, B2 => 
                           n22898, ZN => n4275);
   U14978 : OAI22_X1 port map( A1 => n16646, A2 => n23653, B1 => n19817, B2 => 
                           n22898, ZN => n4281);
   U14979 : OAI22_X1 port map( A1 => n16645, A2 => n23653, B1 => n19816, B2 => 
                           n22898, ZN => n4282);
   U14980 : OAI22_X1 port map( A1 => n16644, A2 => n23653, B1 => n19815, B2 => 
                           n22898, ZN => n4283);
   U14981 : OAI22_X1 port map( A1 => n16643, A2 => n23653, B1 => n19814, B2 => 
                           n22898, ZN => n4284);
   U14982 : OAI22_X1 port map( A1 => n16642, A2 => n23653, B1 => n19813, B2 => 
                           n22898, ZN => n4285);
   U14983 : OAI22_X1 port map( A1 => n16641, A2 => n23653, B1 => n19812, B2 => 
                           n22898, ZN => n4286);
   U14984 : OAI22_X1 port map( A1 => n16640, A2 => n23653, B1 => n19811, B2 => 
                           n22899, ZN => n4287);
   U14985 : OAI22_X1 port map( A1 => n20199, A2 => n23341, B1 => n20263, B2 => 
                           n23333, ZN => n17916);
   U14986 : OAI22_X1 port map( A1 => n19751, A2 => n23398, B1 => n19815, B2 => 
                           n23390, ZN => n17904);
   U14987 : OAI221_X1 port map( B1 => n19943, B2 => n23382, C1 => n19879, C2 =>
                           n23374, A => n17915, ZN => n17903);
   U14988 : AOI222_X1 port map( A1 => n23365, A2 => n21517, B1 => n23357, B2 =>
                           n21088, C1 => n23349, C2 => n20892, ZN => n17915);
   U14989 : OAI22_X1 port map( A1 => n16664, A2 => n23644, B1 => n19899, B2 => 
                           n22891, ZN => n4199);
   U14990 : OAI22_X1 port map( A1 => n16663, A2 => n23643, B1 => n19898, B2 => 
                           n22891, ZN => n4200);
   U14991 : OAI22_X1 port map( A1 => n16662, A2 => n23644, B1 => n19897, B2 => 
                           n22891, ZN => n4201);
   U14992 : OAI22_X1 port map( A1 => n16661, A2 => n23643, B1 => n19896, B2 => 
                           n22891, ZN => n4202);
   U14993 : OAI22_X1 port map( A1 => n16664, A2 => n23664, B1 => n19771, B2 => 
                           n22903, ZN => n4327);
   U14994 : OAI22_X1 port map( A1 => n16663, A2 => n23663, B1 => n19770, B2 => 
                           n22903, ZN => n4328);
   U14995 : OAI22_X1 port map( A1 => n16662, A2 => n23664, B1 => n19769, B2 => 
                           n22903, ZN => n4329);
   U14996 : OAI22_X1 port map( A1 => n16661, A2 => n23663, B1 => n19768, B2 => 
                           n22903, ZN => n4330);
   U14997 : OAI22_X1 port map( A1 => n16664, A2 => n23604, B1 => n20155, B2 => 
                           n22867, ZN => n3943);
   U14998 : OAI22_X1 port map( A1 => n16663, A2 => n23603, B1 => n20154, B2 => 
                           n22867, ZN => n3944);
   U14999 : OAI22_X1 port map( A1 => n16662, A2 => n23604, B1 => n20153, B2 => 
                           n22867, ZN => n3945);
   U15000 : OAI22_X1 port map( A1 => n16661, A2 => n23603, B1 => n20152, B2 => 
                           n22867, ZN => n3946);
   U15001 : OAI22_X1 port map( A1 => n16664, A2 => n23624, B1 => n20027, B2 => 
                           n22879, ZN => n4071);
   U15002 : OAI22_X1 port map( A1 => n16663, A2 => n23623, B1 => n20026, B2 => 
                           n22879, ZN => n4072);
   U15003 : OAI22_X1 port map( A1 => n16662, A2 => n23624, B1 => n20025, B2 => 
                           n22879, ZN => n4073);
   U15004 : OAI22_X1 port map( A1 => n16661, A2 => n23623, B1 => n20024, B2 => 
                           n22879, ZN => n4074);
   U15005 : OAI22_X1 port map( A1 => n16660, A2 => n23654, B1 => n19831, B2 => 
                           n22897, ZN => n4267);
   U15006 : OAI22_X1 port map( A1 => n16659, A2 => n23654, B1 => n19830, B2 => 
                           n22897, ZN => n4268);
   U15007 : OAI22_X1 port map( A1 => n16651, A2 => n23654, B1 => n19822, B2 => 
                           n22898, ZN => n4276);
   U15008 : OAI22_X1 port map( A1 => n16650, A2 => n23654, B1 => n19821, B2 => 
                           n22898, ZN => n4277);
   U15009 : OAI22_X1 port map( A1 => n16649, A2 => n23654, B1 => n19820, B2 => 
                           n22898, ZN => n4278);
   U15010 : OAI22_X1 port map( A1 => n16648, A2 => n23653, B1 => n19819, B2 => 
                           n22898, ZN => n4279);
   U15011 : OAI22_X1 port map( A1 => n16647, A2 => n23653, B1 => n19818, B2 => 
                           n22898, ZN => n4280);
   U15012 : OAI22_X1 port map( A1 => n16639, A2 => n23653, B1 => n19810, B2 => 
                           n22899, ZN => n4288);
   U15013 : OAI22_X1 port map( A1 => n16638, A2 => n23653, B1 => n19809, B2 => 
                           n22899, ZN => n4289);
   U15014 : OAI22_X1 port map( A1 => n16637, A2 => n23653, B1 => n19808, B2 => 
                           n22899, ZN => n4290);
   U15015 : OAI22_X1 port map( A1 => n16658, A2 => n23594, B1 => n20213, B2 => 
                           n22861, ZN => n3885);
   U15016 : OAI22_X1 port map( A1 => n16657, A2 => n23594, B1 => n20212, B2 => 
                           n22861, ZN => n3886);
   U15017 : OAI22_X1 port map( A1 => n16656, A2 => n23594, B1 => n20211, B2 => 
                           n22861, ZN => n3887);
   U15018 : OAI22_X1 port map( A1 => n16655, A2 => n23594, B1 => n20210, B2 => 
                           n22861, ZN => n3888);
   U15019 : OAI22_X1 port map( A1 => n16654, A2 => n23594, B1 => n20209, B2 => 
                           n22861, ZN => n3889);
   U15020 : OAI22_X1 port map( A1 => n16653, A2 => n23594, B1 => n20208, B2 => 
                           n22861, ZN => n3890);
   U15021 : OAI22_X1 port map( A1 => n16652, A2 => n23594, B1 => n20207, B2 => 
                           n22862, ZN => n3891);
   U15022 : OAI22_X1 port map( A1 => n16646, A2 => n23593, B1 => n20201, B2 => 
                           n22862, ZN => n3897);
   U15023 : OAI22_X1 port map( A1 => n16645, A2 => n23593, B1 => n20200, B2 => 
                           n22862, ZN => n3898);
   U15024 : OAI22_X1 port map( A1 => n16644, A2 => n23593, B1 => n20199, B2 => 
                           n22862, ZN => n3899);
   U15025 : OAI22_X1 port map( A1 => n16643, A2 => n23593, B1 => n20198, B2 => 
                           n22862, ZN => n3900);
   U15026 : OAI22_X1 port map( A1 => n16642, A2 => n23593, B1 => n20197, B2 => 
                           n22862, ZN => n3901);
   U15027 : OAI22_X1 port map( A1 => n16641, A2 => n23593, B1 => n20196, B2 => 
                           n22862, ZN => n3902);
   U15028 : OAI22_X1 port map( A1 => n16640, A2 => n23593, B1 => n20195, B2 => 
                           n22863, ZN => n3903);
   U15029 : OAI22_X1 port map( A1 => n16658, A2 => n23614, B1 => n20085, B2 => 
                           n22873, ZN => n4013);
   U15030 : OAI22_X1 port map( A1 => n16657, A2 => n23614, B1 => n20084, B2 => 
                           n22873, ZN => n4014);
   U15031 : OAI22_X1 port map( A1 => n16656, A2 => n23614, B1 => n20083, B2 => 
                           n22873, ZN => n4015);
   U15032 : OAI22_X1 port map( A1 => n16655, A2 => n23614, B1 => n20082, B2 => 
                           n22873, ZN => n4016);
   U15033 : OAI22_X1 port map( A1 => n16654, A2 => n23614, B1 => n20081, B2 => 
                           n22873, ZN => n4017);
   U15034 : OAI22_X1 port map( A1 => n16653, A2 => n23614, B1 => n20080, B2 => 
                           n22873, ZN => n4018);
   U15035 : OAI22_X1 port map( A1 => n16652, A2 => n23614, B1 => n20079, B2 => 
                           n22874, ZN => n4019);
   U15036 : OAI22_X1 port map( A1 => n16646, A2 => n23613, B1 => n20073, B2 => 
                           n22874, ZN => n4025);
   U15037 : OAI22_X1 port map( A1 => n16645, A2 => n23613, B1 => n20072, B2 => 
                           n22874, ZN => n4026);
   U15038 : OAI22_X1 port map( A1 => n16644, A2 => n23613, B1 => n20071, B2 => 
                           n22874, ZN => n4027);
   U15039 : OAI22_X1 port map( A1 => n16643, A2 => n23613, B1 => n20070, B2 => 
                           n22874, ZN => n4028);
   U15040 : OAI22_X1 port map( A1 => n16642, A2 => n23613, B1 => n20069, B2 => 
                           n22874, ZN => n4029);
   U15041 : OAI22_X1 port map( A1 => n16641, A2 => n23613, B1 => n20068, B2 => 
                           n22874, ZN => n4030);
   U15042 : OAI22_X1 port map( A1 => n16640, A2 => n23613, B1 => n20067, B2 => 
                           n22875, ZN => n4031);
   U15043 : OAI22_X1 port map( A1 => n16658, A2 => n23634, B1 => n19957, B2 => 
                           n22885, ZN => n4141);
   U15044 : OAI22_X1 port map( A1 => n16657, A2 => n23634, B1 => n19956, B2 => 
                           n22885, ZN => n4142);
   U15045 : OAI22_X1 port map( A1 => n16656, A2 => n23634, B1 => n19955, B2 => 
                           n22885, ZN => n4143);
   U15046 : OAI22_X1 port map( A1 => n16655, A2 => n23634, B1 => n19954, B2 => 
                           n22885, ZN => n4144);
   U15047 : OAI22_X1 port map( A1 => n16654, A2 => n23634, B1 => n19953, B2 => 
                           n22885, ZN => n4145);
   U15048 : OAI22_X1 port map( A1 => n16653, A2 => n23634, B1 => n19952, B2 => 
                           n22885, ZN => n4146);
   U15049 : OAI22_X1 port map( A1 => n16652, A2 => n23634, B1 => n19951, B2 => 
                           n22886, ZN => n4147);
   U15050 : OAI22_X1 port map( A1 => n16646, A2 => n23633, B1 => n19945, B2 => 
                           n22886, ZN => n4153);
   U15051 : OAI22_X1 port map( A1 => n16645, A2 => n23633, B1 => n19944, B2 => 
                           n22886, ZN => n4154);
   U15052 : OAI22_X1 port map( A1 => n16644, A2 => n23633, B1 => n19943, B2 => 
                           n22886, ZN => n4155);
   U15053 : OAI22_X1 port map( A1 => n16643, A2 => n23633, B1 => n19942, B2 => 
                           n22886, ZN => n4156);
   U15054 : OAI22_X1 port map( A1 => n16642, A2 => n23633, B1 => n19941, B2 => 
                           n22886, ZN => n4157);
   U15055 : OAI22_X1 port map( A1 => n16641, A2 => n23633, B1 => n19940, B2 => 
                           n22886, ZN => n4158);
   U15056 : OAI22_X1 port map( A1 => n16640, A2 => n23633, B1 => n19939, B2 => 
                           n22887, ZN => n4159);
   U15057 : OAI22_X1 port map( A1 => n16660, A2 => n23634, B1 => n19959, B2 => 
                           n22885, ZN => n4139);
   U15058 : OAI22_X1 port map( A1 => n16659, A2 => n23634, B1 => n19958, B2 => 
                           n22885, ZN => n4140);
   U15059 : OAI22_X1 port map( A1 => n16651, A2 => n23634, B1 => n19950, B2 => 
                           n22886, ZN => n4148);
   U15060 : OAI22_X1 port map( A1 => n16650, A2 => n23634, B1 => n19949, B2 => 
                           n22886, ZN => n4149);
   U15061 : OAI22_X1 port map( A1 => n16649, A2 => n23634, B1 => n19948, B2 => 
                           n22886, ZN => n4150);
   U15062 : OAI22_X1 port map( A1 => n16648, A2 => n23633, B1 => n19947, B2 => 
                           n22886, ZN => n4151);
   U15063 : OAI22_X1 port map( A1 => n16647, A2 => n23633, B1 => n19946, B2 => 
                           n22886, ZN => n4152);
   U15064 : OAI22_X1 port map( A1 => n16639, A2 => n23633, B1 => n19938, B2 => 
                           n22887, ZN => n4160);
   U15065 : OAI22_X1 port map( A1 => n16638, A2 => n23633, B1 => n19937, B2 => 
                           n22887, ZN => n4161);
   U15066 : OAI22_X1 port map( A1 => n16637, A2 => n23633, B1 => n19936, B2 => 
                           n22887, ZN => n4162);
   U15067 : OAI22_X1 port map( A1 => n16660, A2 => n23594, B1 => n20215, B2 => 
                           n22861, ZN => n3883);
   U15068 : OAI22_X1 port map( A1 => n16659, A2 => n23594, B1 => n20214, B2 => 
                           n22861, ZN => n3884);
   U15069 : OAI22_X1 port map( A1 => n16651, A2 => n23594, B1 => n20206, B2 => 
                           n22862, ZN => n3892);
   U15070 : OAI22_X1 port map( A1 => n16650, A2 => n23594, B1 => n20205, B2 => 
                           n22862, ZN => n3893);
   U15071 : OAI22_X1 port map( A1 => n16649, A2 => n23594, B1 => n20204, B2 => 
                           n22862, ZN => n3894);
   U15072 : OAI22_X1 port map( A1 => n16648, A2 => n23593, B1 => n20203, B2 => 
                           n22862, ZN => n3895);
   U15073 : OAI22_X1 port map( A1 => n16647, A2 => n23593, B1 => n20202, B2 => 
                           n22862, ZN => n3896);
   U15074 : OAI22_X1 port map( A1 => n16639, A2 => n23593, B1 => n20194, B2 => 
                           n22863, ZN => n3904);
   U15075 : OAI22_X1 port map( A1 => n16638, A2 => n23593, B1 => n20193, B2 => 
                           n22863, ZN => n3905);
   U15076 : OAI22_X1 port map( A1 => n16637, A2 => n23593, B1 => n20192, B2 => 
                           n22863, ZN => n3906);
   U15077 : OAI22_X1 port map( A1 => n16660, A2 => n23614, B1 => n20087, B2 => 
                           n22873, ZN => n4011);
   U15078 : OAI22_X1 port map( A1 => n16659, A2 => n23614, B1 => n20086, B2 => 
                           n22873, ZN => n4012);
   U15079 : OAI22_X1 port map( A1 => n16651, A2 => n23614, B1 => n20078, B2 => 
                           n22874, ZN => n4020);
   U15080 : OAI22_X1 port map( A1 => n16650, A2 => n23614, B1 => n20077, B2 => 
                           n22874, ZN => n4021);
   U15081 : OAI22_X1 port map( A1 => n16649, A2 => n23614, B1 => n20076, B2 => 
                           n22874, ZN => n4022);
   U15082 : OAI22_X1 port map( A1 => n16648, A2 => n23613, B1 => n20075, B2 => 
                           n22874, ZN => n4023);
   U15083 : OAI22_X1 port map( A1 => n16647, A2 => n23613, B1 => n20074, B2 => 
                           n22874, ZN => n4024);
   U15084 : OAI22_X1 port map( A1 => n16639, A2 => n23613, B1 => n20066, B2 => 
                           n22875, ZN => n4032);
   U15085 : OAI22_X1 port map( A1 => n16638, A2 => n23613, B1 => n20065, B2 => 
                           n22875, ZN => n4033);
   U15086 : OAI22_X1 port map( A1 => n16637, A2 => n23613, B1 => n20064, B2 => 
                           n22875, ZN => n4034);
   U15087 : OAI22_X1 port map( A1 => n20187, A2 => n23340, B1 => n20251, B2 => 
                           n23332, ZN => n18483);
   U15088 : OAI22_X1 port map( A1 => n19739, A2 => n23397, B1 => n19803, B2 => 
                           n23389, ZN => n18471);
   U15089 : OAI22_X1 port map( A1 => n20186, A2 => n23340, B1 => n20250, B2 => 
                           n23332, ZN => n18429);
   U15090 : OAI22_X1 port map( A1 => n19738, A2 => n23397, B1 => n19802, B2 => 
                           n23389, ZN => n18417);
   U15091 : OAI22_X1 port map( A1 => n20178, A2 => n23341, B1 => n20242, B2 => 
                           n23333, ZN => n17997);
   U15092 : OAI22_X1 port map( A1 => n19730, A2 => n23398, B1 => n19794, B2 => 
                           n23390, ZN => n17985);
   U15093 : OAI22_X1 port map( A1 => n20193, A2 => n23340, B1 => n20257, B2 => 
                           n23332, ZN => n18240);
   U15094 : OAI22_X1 port map( A1 => n19745, A2 => n23397, B1 => n19809, B2 => 
                           n23389, ZN => n18228);
   U15095 : OAI22_X1 port map( A1 => n20170, A2 => n23342, B1 => n20234, B2 => 
                           n23334, ZN => n17565);
   U15096 : OAI22_X1 port map( A1 => n19722, A2 => n23399, B1 => n19786, B2 => 
                           n23391, ZN => n17553);
   U15097 : OAI22_X1 port map( A1 => n20216, A2 => n23344, B1 => n20280, B2 => 
                           n23336, ZN => n16998);
   U15098 : OAI22_X1 port map( A1 => n19768, A2 => n23401, B1 => n19832, B2 => 
                           n23393, ZN => n16986);
   U15099 : OAI22_X1 port map( A1 => n20179, A2 => n23341, B1 => n20243, B2 => 
                           n23333, ZN => n18051);
   U15100 : OAI22_X1 port map( A1 => n19731, A2 => n23398, B1 => n19795, B2 => 
                           n23390, ZN => n18039);
   U15101 : OAI22_X1 port map( A1 => n20171, A2 => n23342, B1 => n20235, B2 => 
                           n23334, ZN => n17619);
   U15102 : OAI22_X1 port map( A1 => n19723, A2 => n23399, B1 => n19787, B2 => 
                           n23391, ZN => n17607);
   U15103 : OAI22_X1 port map( A1 => n20168, A2 => n23343, B1 => n20232, B2 => 
                           n23335, ZN => n17457);
   U15104 : OAI22_X1 port map( A1 => n19720, A2 => n23400, B1 => n19784, B2 => 
                           n23392, ZN => n17445);
   U15105 : OAI22_X1 port map( A1 => n20167, A2 => n23343, B1 => n20231, B2 => 
                           n23335, ZN => n17403);
   U15106 : OAI22_X1 port map( A1 => n19719, A2 => n23400, B1 => n19783, B2 => 
                           n23392, ZN => n17391);
   U15107 : OAI22_X1 port map( A1 => n20197, A2 => n23341, B1 => n20261, B2 => 
                           n23333, ZN => n18024);
   U15108 : OAI22_X1 port map( A1 => n19749, A2 => n23398, B1 => n19813, B2 => 
                           n23390, ZN => n18012);
   U15109 : OAI22_X1 port map( A1 => n20205, A2 => n23342, B1 => n20269, B2 => 
                           n23334, ZN => n17592);
   U15110 : OAI22_X1 port map( A1 => n19757, A2 => n23399, B1 => n19821, B2 => 
                           n23391, ZN => n17580);
   U15111 : OAI221_X1 port map( B1 => n19931, B2 => n23381, C1 => n19867, C2 =>
                           n23373, A => n18482, ZN => n18470);
   U15112 : AOI222_X1 port map( A1 => n23364, A2 => n21460, B1 => n23356, B2 =>
                           n21031, C1 => n23348, C2 => n20835, ZN => n18482);
   U15113 : OAI221_X1 port map( B1 => n19930, B2 => n23381, C1 => n19866, C2 =>
                           n23373, A => n18428, ZN => n18416);
   U15114 : AOI222_X1 port map( A1 => n23364, A2 => n21475, B1 => n23356, B2 =>
                           n21046, C1 => n23348, C2 => n20850, ZN => n18428);
   U15115 : OAI221_X1 port map( B1 => n19922, B2 => n23382, C1 => n19858, C2 =>
                           n23374, A => n17996, ZN => n17984);
   U15116 : AOI222_X1 port map( A1 => n23365, A2 => n21461, B1 => n23357, B2 =>
                           n21032, C1 => n23349, C2 => n20836, ZN => n17996);
   U15117 : OAI221_X1 port map( B1 => n19937, B2 => n23381, C1 => n19873, C2 =>
                           n23373, A => n18239, ZN => n18227);
   U15118 : AOI222_X1 port map( A1 => n23364, A2 => n21492, B1 => n23356, B2 =>
                           n21063, C1 => n23348, C2 => n20867, ZN => n18239);
   U15119 : OAI221_X1 port map( B1 => n19914, B2 => n23383, C1 => n19850, C2 =>
                           n23375, A => n17564, ZN => n17552);
   U15120 : AOI222_X1 port map( A1 => n23366, A2 => n21462, B1 => n23358, B2 =>
                           n21033, C1 => n23350, C2 => n20837, ZN => n17564);
   U15121 : OAI221_X1 port map( B1 => n19960, B2 => n23385, C1 => n19896, C2 =>
                           n23377, A => n16997, ZN => n16985);
   U15122 : AOI222_X1 port map( A1 => n23368, A2 => n21463, B1 => n23360, B2 =>
                           n21034, C1 => n23352, C2 => n20838, ZN => n16997);
   U15123 : OAI221_X1 port map( B1 => n19923, B2 => n23382, C1 => n19859, C2 =>
                           n23374, A => n18050, ZN => n18038);
   U15124 : AOI222_X1 port map( A1 => n23365, A2 => n21493, B1 => n23357, B2 =>
                           n21064, C1 => n23349, C2 => n20868, ZN => n18050);
   U15125 : OAI221_X1 port map( B1 => n19915, B2 => n23383, C1 => n19851, C2 =>
                           n23375, A => n17618, ZN => n17606);
   U15126 : AOI222_X1 port map( A1 => n23366, A2 => n21464, B1 => n23358, B2 =>
                           n21035, C1 => n23350, C2 => n20839, ZN => n17618);
   U15127 : OAI221_X1 port map( B1 => n19912, B2 => n23384, C1 => n19848, C2 =>
                           n23376, A => n17456, ZN => n17444);
   U15128 : AOI222_X1 port map( A1 => n23367, A2 => n21465, B1 => n23359, B2 =>
                           n21036, C1 => n23351, C2 => n20840, ZN => n17456);
   U15129 : OAI221_X1 port map( B1 => n19911, B2 => n23384, C1 => n19847, C2 =>
                           n23376, A => n17402, ZN => n17390);
   U15130 : AOI222_X1 port map( A1 => n23367, A2 => n21494, B1 => n23359, B2 =>
                           n21065, C1 => n23351, C2 => n20869, ZN => n17402);
   U15131 : OAI221_X1 port map( B1 => n19941, B2 => n23382, C1 => n19877, C2 =>
                           n23374, A => n18023, ZN => n18011);
   U15132 : AOI222_X1 port map( A1 => n23365, A2 => n21476, B1 => n23357, B2 =>
                           n21047, C1 => n23349, C2 => n20851, ZN => n18023);
   U15133 : OAI221_X1 port map( B1 => n19949, B2 => n23383, C1 => n19885, C2 =>
                           n23375, A => n17591, ZN => n17579);
   U15134 : AOI222_X1 port map( A1 => n23366, A2 => n21495, B1 => n23358, B2 =>
                           n21066, C1 => n23350, C2 => n20870, ZN => n17591);
   U15135 : OAI22_X1 port map( A1 => n20194, A2 => n23341, B1 => n20258, B2 => 
                           n23333, ZN => n18186);
   U15136 : OAI22_X1 port map( A1 => n19746, A2 => n23398, B1 => n19810, B2 => 
                           n23390, ZN => n18174);
   U15137 : OAI22_X1 port map( A1 => n20162, A2 => n23344, B1 => n20226, B2 => 
                           n23336, ZN => n17133);
   U15138 : OAI22_X1 port map( A1 => n19714, A2 => n23401, B1 => n19778, B2 => 
                           n23393, ZN => n17121);
   U15139 : OAI22_X1 port map( A1 => n20161, A2 => n23344, B1 => n20225, B2 => 
                           n23336, ZN => n17079);
   U15140 : OAI22_X1 port map( A1 => n19713, A2 => n23401, B1 => n19777, B2 => 
                           n23393, ZN => n17067);
   U15141 : OAI22_X1 port map( A1 => n20160, A2 => n23344, B1 => n20224, B2 => 
                           n23336, ZN => n17025);
   U15142 : OAI22_X1 port map( A1 => n19712, A2 => n23401, B1 => n19776, B2 => 
                           n23393, ZN => n17013);
   U15143 : OAI22_X1 port map( A1 => n20159, A2 => n23344, B1 => n20223, B2 => 
                           n23336, ZN => n16971);
   U15144 : OAI22_X1 port map( A1 => n19711, A2 => n23401, B1 => n19775, B2 => 
                           n23393, ZN => n16959);
   U15145 : OAI22_X1 port map( A1 => n20203, A2 => n23342, B1 => n20267, B2 => 
                           n23334, ZN => n17700);
   U15146 : OAI22_X1 port map( A1 => n19755, A2 => n23399, B1 => n19819, B2 => 
                           n23391, ZN => n17688);
   U15147 : OAI22_X1 port map( A1 => n20210, A2 => n23343, B1 => n20274, B2 => 
                           n23335, ZN => n17322);
   U15148 : OAI22_X1 port map( A1 => n19762, A2 => n23400, B1 => n19826, B2 => 
                           n23392, ZN => n17310);
   U15149 : OAI22_X1 port map( A1 => n20190, A2 => n23340, B1 => n20254, B2 => 
                           n23332, ZN => n18402);
   U15150 : OAI22_X1 port map( A1 => n19742, A2 => n23397, B1 => n19806, B2 => 
                           n23389, ZN => n18390);
   U15151 : OAI22_X1 port map( A1 => n20191, A2 => n23340, B1 => n20255, B2 => 
                           n23332, ZN => n18348);
   U15152 : OAI22_X1 port map( A1 => n19743, A2 => n23397, B1 => n19807, B2 => 
                           n23389, ZN => n18336);
   U15153 : OAI22_X1 port map( A1 => n20176, A2 => n23341, B1 => n20240, B2 => 
                           n23333, ZN => n17889);
   U15154 : OAI22_X1 port map( A1 => n19728, A2 => n23398, B1 => n19792, B2 => 
                           n23390, ZN => n17877);
   U15155 : OAI22_X1 port map( A1 => n20173, A2 => n23342, B1 => n20237, B2 => 
                           n23334, ZN => n17727);
   U15156 : OAI22_X1 port map( A1 => n19725, A2 => n23399, B1 => n19789, B2 => 
                           n23391, ZN => n17715);
   U15157 : OAI22_X1 port map( A1 => n20172, A2 => n23342, B1 => n20236, B2 => 
                           n23334, ZN => n17673);
   U15158 : OAI22_X1 port map( A1 => n19724, A2 => n23399, B1 => n19788, B2 => 
                           n23391, ZN => n17661);
   U15159 : OAI22_X1 port map( A1 => n20207, A2 => n23343, B1 => n20271, B2 => 
                           n23335, ZN => n17484);
   U15160 : OAI22_X1 port map( A1 => n19759, A2 => n23400, B1 => n19823, B2 => 
                           n23392, ZN => n17472);
   U15161 : OAI22_X1 port map( A1 => n20164, A2 => n23343, B1 => n20228, B2 => 
                           n23335, ZN => n17241);
   U15162 : OAI22_X1 port map( A1 => n19716, A2 => n23400, B1 => n19780, B2 => 
                           n23392, ZN => n17229);
   U15163 : OAI22_X1 port map( A1 => n20215, A2 => n23344, B1 => n20279, B2 => 
                           n23336, ZN => n17052);
   U15164 : OAI22_X1 port map( A1 => n19767, A2 => n23401, B1 => n19831, B2 => 
                           n23393, ZN => n17040);
   U15165 : OAI22_X1 port map( A1 => n20182, A2 => n23340, B1 => n20246, B2 => 
                           n23332, ZN => n18213);
   U15166 : OAI22_X1 port map( A1 => n19734, A2 => n23397, B1 => n19798, B2 => 
                           n23389, ZN => n18201);
   U15167 : OAI22_X1 port map( A1 => n20195, A2 => n23341, B1 => n20259, B2 => 
                           n23333, ZN => n18132);
   U15168 : OAI22_X1 port map( A1 => n19747, A2 => n23398, B1 => n19811, B2 => 
                           n23390, ZN => n18120);
   U15169 : OAI22_X1 port map( A1 => n20204, A2 => n23342, B1 => n20268, B2 => 
                           n23334, ZN => n17646);
   U15170 : OAI22_X1 port map( A1 => n19756, A2 => n23399, B1 => n19820, B2 => 
                           n23391, ZN => n17634);
   U15171 : OAI22_X1 port map( A1 => n20196, A2 => n23341, B1 => n20260, B2 => 
                           n23333, ZN => n18078);
   U15172 : OAI22_X1 port map( A1 => n19748, A2 => n23398, B1 => n19812, B2 => 
                           n23390, ZN => n18066);
   U15173 : OAI22_X1 port map( A1 => n20198, A2 => n23341, B1 => n20262, B2 => 
                           n23333, ZN => n17970);
   U15174 : OAI22_X1 port map( A1 => n19750, A2 => n23398, B1 => n19814, B2 => 
                           n23390, ZN => n17958);
   U15175 : OAI22_X1 port map( A1 => n20209, A2 => n23343, B1 => n20273, B2 => 
                           n23335, ZN => n17376);
   U15176 : OAI22_X1 port map( A1 => n19761, A2 => n23400, B1 => n19825, B2 => 
                           n23392, ZN => n17364);
   U15177 : OAI22_X1 port map( A1 => n20165, A2 => n23343, B1 => n20229, B2 => 
                           n23335, ZN => n17295);
   U15178 : OAI22_X1 port map( A1 => n19717, A2 => n23400, B1 => n19781, B2 => 
                           n23392, ZN => n17283);
   U15179 : OAI22_X1 port map( A1 => n20163, A2 => n23344, B1 => n20227, B2 => 
                           n23336, ZN => n17187);
   U15180 : OAI22_X1 port map( A1 => n19715, A2 => n23401, B1 => n19779, B2 => 
                           n23393, ZN => n17175);
   U15181 : OAI22_X1 port map( A1 => n20217, A2 => n23344, B1 => n20281, B2 => 
                           n23336, ZN => n16944);
   U15182 : OAI22_X1 port map( A1 => n19769, A2 => n23401, B1 => n19833, B2 => 
                           n23393, ZN => n16932);
   U15183 : OAI22_X1 port map( A1 => n20189, A2 => n23340, B1 => n20253, B2 => 
                           n23332, ZN => n18456);
   U15184 : OAI22_X1 port map( A1 => n19741, A2 => n23397, B1 => n19805, B2 => 
                           n23389, ZN => n18444);
   U15185 : OAI22_X1 port map( A1 => n20183, A2 => n23340, B1 => n20247, B2 => 
                           n23332, ZN => n18267);
   U15186 : OAI22_X1 port map( A1 => n19735, A2 => n23397, B1 => n19799, B2 => 
                           n23389, ZN => n18255);
   U15187 : OAI22_X1 port map( A1 => n20174, A2 => n23342, B1 => n20238, B2 => 
                           n23334, ZN => n17781);
   U15188 : OAI22_X1 port map( A1 => n19726, A2 => n23399, B1 => n19790, B2 => 
                           n23391, ZN => n17769);
   U15189 : OAI22_X1 port map( A1 => n20166, A2 => n23343, B1 => n20230, B2 => 
                           n23335, ZN => n17349);
   U15190 : OAI22_X1 port map( A1 => n19718, A2 => n23400, B1 => n19782, B2 => 
                           n23392, ZN => n17337);
   U15191 : OAI22_X1 port map( A1 => n20211, A2 => n23343, B1 => n20275, B2 => 
                           n23335, ZN => n17268);
   U15192 : OAI22_X1 port map( A1 => n19763, A2 => n23400, B1 => n19827, B2 => 
                           n23392, ZN => n17256);
   U15193 : OAI22_X1 port map( A1 => n20212, A2 => n23344, B1 => n20276, B2 => 
                           n23336, ZN => n17214);
   U15194 : OAI22_X1 port map( A1 => n19764, A2 => n23401, B1 => n19828, B2 => 
                           n23393, ZN => n17202);
   U15195 : OAI22_X1 port map( A1 => n20213, A2 => n23344, B1 => n20277, B2 => 
                           n23336, ZN => n17160);
   U15196 : OAI22_X1 port map( A1 => n19765, A2 => n23401, B1 => n19829, B2 => 
                           n23393, ZN => n17148);
   U15197 : OAI22_X1 port map( A1 => n20214, A2 => n23344, B1 => n20278, B2 => 
                           n23336, ZN => n17106);
   U15198 : OAI22_X1 port map( A1 => n19766, A2 => n23401, B1 => n19830, B2 => 
                           n23393, ZN => n17094);
   U15199 : OAI22_X1 port map( A1 => n20158, A2 => n23344, B1 => n20222, B2 => 
                           n23336, ZN => n16917);
   U15200 : OAI22_X1 port map( A1 => n19710, A2 => n23401, B1 => n19774, B2 => 
                           n23393, ZN => n16905);
   U15201 : OAI22_X1 port map( A1 => n20206, A2 => n23343, B1 => n20270, B2 => 
                           n23335, ZN => n17538);
   U15202 : OAI22_X1 port map( A1 => n19758, A2 => n23400, B1 => n19822, B2 => 
                           n23392, ZN => n17526);
   U15203 : OAI22_X1 port map( A1 => n20208, A2 => n23343, B1 => n20272, B2 => 
                           n23335, ZN => n17430);
   U15204 : OAI22_X1 port map( A1 => n19760, A2 => n23400, B1 => n19824, B2 => 
                           n23392, ZN => n17418);
   U15205 : OAI221_X1 port map( B1 => n19938, B2 => n23382, C1 => n19874, C2 =>
                           n23374, A => n18185, ZN => n18173);
   U15206 : AOI222_X1 port map( A1 => n23365, A2 => n21477, B1 => n23357, B2 =>
                           n21048, C1 => n23349, C2 => n20852, ZN => n18185);
   U15207 : OAI221_X1 port map( B1 => n19906, B2 => n23385, C1 => n19842, C2 =>
                           n23377, A => n17132, ZN => n17120);
   U15208 : AOI222_X1 port map( A1 => n23368, A2 => n21496, B1 => n23360, B2 =>
                           n21067, C1 => n23352, C2 => n20871, ZN => n17132);
   U15209 : OAI221_X1 port map( B1 => n19905, B2 => n23385, C1 => n19841, C2 =>
                           n23377, A => n17078, ZN => n17066);
   U15210 : AOI222_X1 port map( A1 => n23368, A2 => n21466, B1 => n23360, B2 =>
                           n21037, C1 => n23352, C2 => n20841, ZN => n17078);
   U15211 : OAI221_X1 port map( B1 => n19904, B2 => n23385, C1 => n19840, C2 =>
                           n23377, A => n17024, ZN => n17012);
   U15212 : AOI222_X1 port map( A1 => n23368, A2 => n21497, B1 => n23360, B2 =>
                           n21068, C1 => n23352, C2 => n20872, ZN => n17024);
   U15213 : OAI221_X1 port map( B1 => n19903, B2 => n23385, C1 => n19839, C2 =>
                           n23377, A => n16970, ZN => n16958);
   U15214 : AOI222_X1 port map( A1 => n23368, A2 => n21498, B1 => n23360, B2 =>
                           n21069, C1 => n23352, C2 => n20873, ZN => n16970);
   U15215 : OAI221_X1 port map( B1 => n19947, B2 => n23383, C1 => n19883, C2 =>
                           n23375, A => n17699, ZN => n17687);
   U15216 : AOI222_X1 port map( A1 => n23366, A2 => n21478, B1 => n23358, B2 =>
                           n21049, C1 => n23350, C2 => n20853, ZN => n17699);
   U15217 : OAI221_X1 port map( B1 => n19954, B2 => n23384, C1 => n19890, C2 =>
                           n23376, A => n17321, ZN => n17309);
   U15218 : AOI222_X1 port map( A1 => n23367, A2 => n21467, B1 => n23359, B2 =>
                           n21038, C1 => n23351, C2 => n20842, ZN => n17321);
   U15219 : OAI221_X1 port map( B1 => n19934, B2 => n23381, C1 => n19870, C2 =>
                           n23373, A => n18401, ZN => n18389);
   U15220 : AOI222_X1 port map( A1 => n23364, A2 => n21479, B1 => n23356, B2 =>
                           n21050, C1 => n23348, C2 => n20854, ZN => n18401);
   U15221 : OAI221_X1 port map( B1 => n19935, B2 => n23381, C1 => n19871, C2 =>
                           n23373, A => n18347, ZN => n18335);
   U15222 : AOI222_X1 port map( A1 => n23364, A2 => n21480, B1 => n23356, B2 =>
                           n21051, C1 => n23348, C2 => n20855, ZN => n18347);
   U15223 : OAI221_X1 port map( B1 => n19920, B2 => n23382, C1 => n19856, C2 =>
                           n23374, A => n17888, ZN => n17876);
   U15224 : AOI222_X1 port map( A1 => n23365, A2 => n21481, B1 => n23357, B2 =>
                           n21052, C1 => n23349, C2 => n20856, ZN => n17888);
   U15225 : OAI221_X1 port map( B1 => n19917, B2 => n23383, C1 => n19853, C2 =>
                           n23375, A => n17726, ZN => n17714);
   U15226 : AOI222_X1 port map( A1 => n23366, A2 => n21482, B1 => n23358, B2 =>
                           n21053, C1 => n23350, C2 => n20857, ZN => n17726);
   U15227 : OAI221_X1 port map( B1 => n19916, B2 => n23383, C1 => n19852, C2 =>
                           n23375, A => n17672, ZN => n17660);
   U15228 : AOI222_X1 port map( A1 => n23366, A2 => n21483, B1 => n23358, B2 =>
                           n21054, C1 => n23350, C2 => n20858, ZN => n17672);
   U15229 : OAI221_X1 port map( B1 => n19951, B2 => n23384, C1 => n19887, C2 =>
                           n23376, A => n17483, ZN => n17471);
   U15230 : AOI222_X1 port map( A1 => n23367, A2 => n21484, B1 => n23359, B2 =>
                           n21055, C1 => n23351, C2 => n20859, ZN => n17483);
   U15231 : OAI221_X1 port map( B1 => n19908, B2 => n23384, C1 => n19844, C2 =>
                           n23376, A => n17240, ZN => n17228);
   U15232 : AOI222_X1 port map( A1 => n23367, A2 => n21468, B1 => n23359, B2 =>
                           n21039, C1 => n23351, C2 => n20843, ZN => n17240);
   U15233 : OAI221_X1 port map( B1 => n19959, B2 => n23385, C1 => n19895, C2 =>
                           n23377, A => n17051, ZN => n17039);
   U15234 : AOI222_X1 port map( A1 => n23368, A2 => n21499, B1 => n23360, B2 =>
                           n21070, C1 => n23352, C2 => n20874, ZN => n17051);
   U15235 : OAI221_X1 port map( B1 => n19926, B2 => n23381, C1 => n19862, C2 =>
                           n23373, A => n18212, ZN => n18200);
   U15236 : AOI222_X1 port map( A1 => n23364, A2 => n21485, B1 => n23356, B2 =>
                           n21056, C1 => n23348, C2 => n20860, ZN => n18212);
   U15237 : OAI221_X1 port map( B1 => n19939, B2 => n23382, C1 => n19875, C2 =>
                           n23374, A => n18131, ZN => n18119);
   U15238 : AOI222_X1 port map( A1 => n23365, A2 => n21486, B1 => n23357, B2 =>
                           n21057, C1 => n23349, C2 => n20861, ZN => n18131);
   U15239 : OAI221_X1 port map( B1 => n19948, B2 => n23383, C1 => n19884, C2 =>
                           n23375, A => n17645, ZN => n17633);
   U15240 : AOI222_X1 port map( A1 => n23366, A2 => n21520, B1 => n23358, B2 =>
                           n21091, C1 => n23350, C2 => n20895, ZN => n17645);
   U15241 : OAI221_X1 port map( B1 => n19940, B2 => n23382, C1 => n19876, C2 =>
                           n23374, A => n18077, ZN => n18065);
   U15242 : AOI222_X1 port map( A1 => n23365, A2 => n21487, B1 => n23357, B2 =>
                           n21058, C1 => n23349, C2 => n20862, ZN => n18077);
   U15243 : OAI221_X1 port map( B1 => n19942, B2 => n23382, C1 => n19878, C2 =>
                           n23374, A => n17969, ZN => n17957);
   U15244 : AOI222_X1 port map( A1 => n23365, A2 => n21488, B1 => n23357, B2 =>
                           n21059, C1 => n23349, C2 => n20863, ZN => n17969);
   U15245 : OAI221_X1 port map( B1 => n19953, B2 => n23384, C1 => n19889, C2 =>
                           n23376, A => n17375, ZN => n17363);
   U15246 : AOI222_X1 port map( A1 => n23367, A2 => n21469, B1 => n23359, B2 =>
                           n21040, C1 => n23351, C2 => n20844, ZN => n17375);
   U15247 : OAI221_X1 port map( B1 => n19909, B2 => n23384, C1 => n19845, C2 =>
                           n23376, A => n17294, ZN => n17282);
   U15248 : AOI222_X1 port map( A1 => n23367, A2 => n21500, B1 => n23359, B2 =>
                           n21071, C1 => n23351, C2 => n20875, ZN => n17294);
   U15249 : OAI221_X1 port map( B1 => n19907, B2 => n23385, C1 => n19843, C2 =>
                           n23377, A => n17186, ZN => n17174);
   U15250 : AOI222_X1 port map( A1 => n23368, A2 => n21489, B1 => n23360, B2 =>
                           n21060, C1 => n23352, C2 => n20864, ZN => n17186);
   U15251 : OAI221_X1 port map( B1 => n19961, B2 => n23385, C1 => n19897, C2 =>
                           n23377, A => n16943, ZN => n16931);
   U15252 : AOI222_X1 port map( A1 => n23368, A2 => n21501, B1 => n23360, B2 =>
                           n21072, C1 => n23352, C2 => n20876, ZN => n16943);
   U15253 : OAI221_X1 port map( B1 => n19933, B2 => n23381, C1 => n19869, C2 =>
                           n23373, A => n18455, ZN => n18443);
   U15254 : AOI222_X1 port map( A1 => n23364, A2 => n21490, B1 => n23356, B2 =>
                           n21061, C1 => n23348, C2 => n20865, ZN => n18455);
   U15255 : OAI221_X1 port map( B1 => n19927, B2 => n23381, C1 => n19863, C2 =>
                           n23373, A => n18266, ZN => n18254);
   U15256 : AOI222_X1 port map( A1 => n23364, A2 => n21516, B1 => n23356, B2 =>
                           n21087, C1 => n23348, C2 => n20891, ZN => n18266);
   U15257 : OAI221_X1 port map( B1 => n19918, B2 => n23383, C1 => n19854, C2 =>
                           n23375, A => n17780, ZN => n17768);
   U15258 : AOI222_X1 port map( A1 => n23366, A2 => n21491, B1 => n23358, B2 =>
                           n21062, C1 => n23350, C2 => n20866, ZN => n17780);
   U15259 : OAI221_X1 port map( B1 => n19910, B2 => n23384, C1 => n19846, C2 =>
                           n23376, A => n17348, ZN => n17336);
   U15260 : AOI222_X1 port map( A1 => n23367, A2 => n21502, B1 => n23359, B2 =>
                           n21073, C1 => n23351, C2 => n20877, ZN => n17348);
   U15261 : OAI221_X1 port map( B1 => n19955, B2 => n23384, C1 => n19891, C2 =>
                           n23376, A => n17267, ZN => n17255);
   U15262 : AOI222_X1 port map( A1 => n23367, A2 => n21503, B1 => n23359, B2 =>
                           n21074, C1 => n23351, C2 => n20878, ZN => n17267);
   U15263 : OAI221_X1 port map( B1 => n19956, B2 => n23385, C1 => n19892, C2 =>
                           n23377, A => n17213, ZN => n17201);
   U15264 : AOI222_X1 port map( A1 => n23368, A2 => n21504, B1 => n23360, B2 =>
                           n21075, C1 => n23352, C2 => n20879, ZN => n17213);
   U15265 : OAI221_X1 port map( B1 => n19957, B2 => n23385, C1 => n19893, C2 =>
                           n23377, A => n17159, ZN => n17147);
   U15266 : AOI222_X1 port map( A1 => n23368, A2 => n21470, B1 => n23360, B2 =>
                           n21041, C1 => n23352, C2 => n20845, ZN => n17159);
   U15267 : OAI221_X1 port map( B1 => n19958, B2 => n23385, C1 => n19894, C2 =>
                           n23377, A => n17105, ZN => n17093);
   U15268 : AOI222_X1 port map( A1 => n23368, A2 => n21505, B1 => n23360, B2 =>
                           n21076, C1 => n23352, C2 => n20880, ZN => n17105);
   U15269 : OAI221_X1 port map( B1 => n19902, B2 => n23385, C1 => n19838, C2 =>
                           n23377, A => n16916, ZN => n16904);
   U15270 : AOI222_X1 port map( A1 => n23368, A2 => n21471, B1 => n23360, B2 =>
                           n21042, C1 => n23352, C2 => n20846, ZN => n16916);
   U15271 : OAI221_X1 port map( B1 => n19950, B2 => n23384, C1 => n19886, C2 =>
                           n23376, A => n17537, ZN => n17525);
   U15272 : AOI222_X1 port map( A1 => n23367, A2 => n21521, B1 => n23359, B2 =>
                           n21092, C1 => n23351, C2 => n20896, ZN => n17537);
   U15273 : OAI221_X1 port map( B1 => n19952, B2 => n23384, C1 => n19888, C2 =>
                           n23376, A => n17429, ZN => n17417);
   U15274 : AOI222_X1 port map( A1 => n23367, A2 => n21518, B1 => n23359, B2 =>
                           n21089, C1 => n23351, C2 => n20893, ZN => n17429);
   U15275 : OAI22_X1 port map( A1 => n16664, A2 => n23654, B1 => n19835, B2 => 
                           n22897, ZN => n4263);
   U15276 : OAI22_X1 port map( A1 => n16663, A2 => n23653, B1 => n19834, B2 => 
                           n22897, ZN => n4264);
   U15277 : OAI22_X1 port map( A1 => n16662, A2 => n23654, B1 => n19833, B2 => 
                           n22897, ZN => n4265);
   U15278 : OAI22_X1 port map( A1 => n16661, A2 => n23653, B1 => n19832, B2 => 
                           n22897, ZN => n4266);
   U15279 : OAI22_X1 port map( A1 => n20192, A2 => n23340, B1 => n20256, B2 => 
                           n23332, ZN => n18294);
   U15280 : OAI22_X1 port map( A1 => n19744, A2 => n23397, B1 => n19808, B2 => 
                           n23389, ZN => n18282);
   U15281 : OAI22_X1 port map( A1 => n20200, A2 => n23342, B1 => n20264, B2 => 
                           n23334, ZN => n17862);
   U15282 : OAI22_X1 port map( A1 => n19752, A2 => n23399, B1 => n19816, B2 => 
                           n23391, ZN => n17850);
   U15283 : OAI221_X1 port map( B1 => n19936, B2 => n23381, C1 => n19872, C2 =>
                           n23373, A => n18293, ZN => n18281);
   U15284 : AOI222_X1 port map( A1 => n23364, A2 => n21506, B1 => n23356, B2 =>
                           n21077, C1 => n23348, C2 => n20881, ZN => n18293);
   U15285 : OAI221_X1 port map( B1 => n19944, B2 => n23383, C1 => n19880, C2 =>
                           n23375, A => n17861, ZN => n17849);
   U15286 : AOI222_X1 port map( A1 => n23366, A2 => n21472, B1 => n23358, B2 =>
                           n21043, C1 => n23350, C2 => n20847, ZN => n17861);
   U15287 : OAI22_X1 port map( A1 => n20185, A2 => n23340, B1 => n20249, B2 => 
                           n23332, ZN => n18375);
   U15288 : OAI22_X1 port map( A1 => n19737, A2 => n23397, B1 => n19801, B2 => 
                           n23389, ZN => n18363);
   U15289 : OAI22_X1 port map( A1 => n20201, A2 => n23342, B1 => n20265, B2 => 
                           n23334, ZN => n17808);
   U15290 : OAI22_X1 port map( A1 => n19753, A2 => n23399, B1 => n19817, B2 => 
                           n23391, ZN => n17796);
   U15291 : OAI22_X1 port map( A1 => n20202, A2 => n23342, B1 => n20266, B2 => 
                           n23334, ZN => n17754);
   U15292 : OAI22_X1 port map( A1 => n19754, A2 => n23399, B1 => n19818, B2 => 
                           n23391, ZN => n17742);
   U15293 : OAI22_X1 port map( A1 => n20184, A2 => n23340, B1 => n20248, B2 => 
                           n23332, ZN => n18321);
   U15294 : OAI22_X1 port map( A1 => n19736, A2 => n23397, B1 => n19800, B2 => 
                           n23389, ZN => n18309);
   U15295 : OAI22_X1 port map( A1 => n20181, A2 => n23341, B1 => n20245, B2 => 
                           n23333, ZN => n18159);
   U15296 : OAI22_X1 port map( A1 => n19733, A2 => n23398, B1 => n19797, B2 => 
                           n23390, ZN => n18147);
   U15297 : OAI22_X1 port map( A1 => n20180, A2 => n23341, B1 => n20244, B2 => 
                           n23333, ZN => n18105);
   U15298 : OAI22_X1 port map( A1 => n19732, A2 => n23398, B1 => n19796, B2 => 
                           n23390, ZN => n18093);
   U15299 : OAI22_X1 port map( A1 => n20177, A2 => n23341, B1 => n20241, B2 => 
                           n23333, ZN => n17943);
   U15300 : OAI22_X1 port map( A1 => n19729, A2 => n23398, B1 => n19793, B2 => 
                           n23390, ZN => n17931);
   U15301 : OAI22_X1 port map( A1 => n20175, A2 => n23342, B1 => n20239, B2 => 
                           n23334, ZN => n17835);
   U15302 : OAI22_X1 port map( A1 => n19727, A2 => n23399, B1 => n19791, B2 => 
                           n23391, ZN => n17823);
   U15303 : OAI221_X1 port map( B1 => n19929, B2 => n23381, C1 => n19865, C2 =>
                           n23373, A => n18374, ZN => n18362);
   U15304 : AOI222_X1 port map( A1 => n23364, A2 => n21473, B1 => n23356, B2 =>
                           n21044, C1 => n23348, C2 => n20848, ZN => n18374);
   U15305 : OAI221_X1 port map( B1 => n19945, B2 => n23383, C1 => n19881, C2 =>
                           n23375, A => n17807, ZN => n17795);
   U15306 : AOI222_X1 port map( A1 => n23366, A2 => n21474, B1 => n23358, B2 =>
                           n21045, C1 => n23350, C2 => n20849, ZN => n17807);
   U15307 : OAI221_X1 port map( B1 => n19946, B2 => n23383, C1 => n19882, C2 =>
                           n23375, A => n17753, ZN => n17741);
   U15308 : AOI222_X1 port map( A1 => n23366, A2 => n21507, B1 => n23358, B2 =>
                           n21078, C1 => n23350, C2 => n20882, ZN => n17753);
   U15309 : OAI221_X1 port map( B1 => n19928, B2 => n23381, C1 => n19864, C2 =>
                           n23373, A => n18320, ZN => n18308);
   U15310 : AOI222_X1 port map( A1 => n23364, A2 => n21508, B1 => n23356, B2 =>
                           n21079, C1 => n23348, C2 => n20883, ZN => n18320);
   U15311 : OAI221_X1 port map( B1 => n19925, B2 => n23382, C1 => n19861, C2 =>
                           n23374, A => n18158, ZN => n18146);
   U15312 : AOI222_X1 port map( A1 => n23365, A2 => n21509, B1 => n23357, B2 =>
                           n21080, C1 => n23349, C2 => n20884, ZN => n18158);
   U15313 : OAI221_X1 port map( B1 => n19924, B2 => n23382, C1 => n19860, C2 =>
                           n23374, A => n18104, ZN => n18092);
   U15314 : AOI222_X1 port map( A1 => n23365, A2 => n21519, B1 => n23357, B2 =>
                           n21090, C1 => n23349, C2 => n20894, ZN => n18104);
   U15315 : OAI221_X1 port map( B1 => n19921, B2 => n23382, C1 => n19857, C2 =>
                           n23374, A => n17942, ZN => n17930);
   U15316 : AOI222_X1 port map( A1 => n23365, A2 => n21510, B1 => n23357, B2 =>
                           n21081, C1 => n23349, C2 => n20885, ZN => n17942);
   U15317 : OAI221_X1 port map( B1 => n19919, B2 => n23383, C1 => n19855, C2 =>
                           n23375, A => n17834, ZN => n17822);
   U15318 : AOI222_X1 port map( A1 => n23366, A2 => n21511, B1 => n23358, B2 =>
                           n21082, C1 => n23350, C2 => n20886, ZN => n17834);
   U15319 : OAI22_X1 port map( A1 => n16664, A2 => n23634, B1 => n19963, B2 => 
                           n22885, ZN => n4135);
   U15320 : OAI22_X1 port map( A1 => n16663, A2 => n23633, B1 => n19962, B2 => 
                           n22885, ZN => n4136);
   U15321 : OAI22_X1 port map( A1 => n16662, A2 => n23634, B1 => n19961, B2 => 
                           n22885, ZN => n4137);
   U15322 : OAI22_X1 port map( A1 => n16661, A2 => n23633, B1 => n19960, B2 => 
                           n22885, ZN => n4138);
   U15323 : OAI22_X1 port map( A1 => n16664, A2 => n23594, B1 => n20219, B2 => 
                           n22861, ZN => n3879);
   U15324 : OAI22_X1 port map( A1 => n16663, A2 => n23593, B1 => n20218, B2 => 
                           n22861, ZN => n3880);
   U15325 : OAI22_X1 port map( A1 => n16662, A2 => n23594, B1 => n20217, B2 => 
                           n22861, ZN => n3881);
   U15326 : OAI22_X1 port map( A1 => n16661, A2 => n23593, B1 => n20216, B2 => 
                           n22861, ZN => n3882);
   U15327 : OAI22_X1 port map( A1 => n16664, A2 => n23614, B1 => n20091, B2 => 
                           n22873, ZN => n4007);
   U15328 : OAI22_X1 port map( A1 => n16663, A2 => n23613, B1 => n20090, B2 => 
                           n22873, ZN => n4008);
   U15329 : OAI22_X1 port map( A1 => n16662, A2 => n23614, B1 => n20089, B2 => 
                           n22873, ZN => n4009);
   U15330 : OAI22_X1 port map( A1 => n16661, A2 => n23613, B1 => n20088, B2 => 
                           n22873, ZN => n4010);
   U15331 : OAI22_X1 port map( A1 => n20218, A2 => n23345, B1 => n20282, B2 => 
                           n23337, ZN => n16890);
   U15332 : OAI22_X1 port map( A1 => n19770, A2 => n23402, B1 => n19834, B2 => 
                           n23394, ZN => n16878);
   U15333 : OAI22_X1 port map( A1 => n20219, A2 => n23345, B1 => n20283, B2 => 
                           n23337, ZN => n16836);
   U15334 : OAI22_X1 port map( A1 => n19771, A2 => n23402, B1 => n19835, B2 => 
                           n23394, ZN => n16824);
   U15335 : OAI221_X1 port map( B1 => n19962, B2 => n23386, C1 => n19898, C2 =>
                           n23378, A => n16889, ZN => n16877);
   U15336 : AOI222_X1 port map( A1 => n23369, A2 => n21513, B1 => n23361, B2 =>
                           n21084, C1 => n23353, C2 => n20888, ZN => n16889);
   U15337 : OAI221_X1 port map( B1 => n19963, B2 => n23386, C1 => n19899, C2 =>
                           n23378, A => n16835, ZN => n16823);
   U15338 : AOI222_X1 port map( A1 => n23369, A2 => n21512, B1 => n23361, B2 =>
                           n21083, C1 => n23353, C2 => n20887, ZN => n16835);
   U15339 : OAI22_X1 port map( A1 => n20157, A2 => n23345, B1 => n20221, B2 => 
                           n23337, ZN => n16863);
   U15340 : OAI22_X1 port map( A1 => n19709, A2 => n23402, B1 => n19773, B2 => 
                           n23394, ZN => n16851);
   U15341 : OAI22_X1 port map( A1 => n20156, A2 => n23345, B1 => n20220, B2 => 
                           n23337, ZN => n16802);
   U15342 : OAI22_X1 port map( A1 => n19708, A2 => n23402, B1 => n19772, B2 => 
                           n23394, ZN => n16771);
   U15343 : OAI221_X1 port map( B1 => n19901, B2 => n23386, C1 => n19837, C2 =>
                           n23378, A => n16862, ZN => n16850);
   U15344 : AOI222_X1 port map( A1 => n23369, A2 => n21514, B1 => n23361, B2 =>
                           n21085, C1 => n23353, C2 => n20889, ZN => n16862);
   U15345 : OAI221_X1 port map( B1 => n19900, B2 => n23386, C1 => n19836, C2 =>
                           n23378, A => n16796, ZN => n16770);
   U15346 : AOI222_X1 port map( A1 => n23369, A2 => n21515, B1 => n23361, B2 =>
                           n21086, C1 => n23353, C2 => n20890, ZN => n16796);
   U15347 : OAI221_X1 port map( B1 => n19913, B2 => n23384, C1 => n19849, C2 =>
                           n23376, A => n17510, ZN => n17498);
   U15348 : AOI222_X1 port map( A1 => n23367, A2 => n21522, B1 => n23359, B2 =>
                           n21093, C1 => n23351, C2 => n20897, ZN => n17510);
   U15349 : OAI221_X1 port map( B1 => n19932, B2 => n23381, C1 => n19868, C2 =>
                           n23373, A => n18522, ZN => n18509);
   U15350 : AOI222_X1 port map( A1 => n23364, A2 => n21763, B1 => n23356, B2 =>
                           n21272, C1 => n23348, C2 => n20898, ZN => n18522);
   U15351 : OAI22_X1 port map( A1 => n19721, A2 => n23400, B1 => n19785, B2 => 
                           n23392, ZN => n17499);
   U15352 : OAI22_X1 port map( A1 => n20169, A2 => n23343, B1 => n20233, B2 => 
                           n23335, ZN => n17511);
   U15353 : OAI22_X1 port map( A1 => n19740, A2 => n23397, B1 => n19804, B2 => 
                           n23389, ZN => n18510);
   U15354 : OAI22_X1 port map( A1 => n20188, A2 => n23340, B1 => n20252, B2 => 
                           n23332, ZN => n18523);
   U15355 : BUF_X1 port map( A => n15181, Z => n23908);
   U15356 : OAI22_X1 port map( A1 => n18780, A2 => n23918, B1 => n18844, B2 => 
                           n23909, ZN => n16528);
   U15357 : AND2_X1 port map( A1 => n23283, A2 => n16581, ZN => n22766);
   U15358 : OAI22_X1 port map( A1 => n18748, A2 => n23918, B1 => n18812, B2 => 
                           n23909, ZN => n16507);
   U15359 : OAI22_X1 port map( A1 => n18811, A2 => n23918, B1 => n18875, B2 => 
                           n23909, ZN => n16486);
   U15360 : OAI22_X1 port map( A1 => n18749, A2 => n23918, B1 => n18813, B2 => 
                           n23909, ZN => n16465);
   U15361 : OAI22_X1 port map( A1 => n18810, A2 => n23918, B1 => n18874, B2 => 
                           n23909, ZN => n16444);
   U15362 : OAI22_X1 port map( A1 => n18750, A2 => n23918, B1 => n18814, B2 => 
                           n23909, ZN => n16423);
   U15363 : OAI22_X1 port map( A1 => n18809, A2 => n23918, B1 => n18873, B2 => 
                           n23909, ZN => n16402);
   U15364 : OAI22_X1 port map( A1 => n18751, A2 => n23918, B1 => n18815, B2 => 
                           n23909, ZN => n16381);
   U15365 : OAI22_X1 port map( A1 => n18808, A2 => n23918, B1 => n18872, B2 => 
                           n23909, ZN => n16360);
   U15366 : OAI22_X1 port map( A1 => n18752, A2 => n23918, B1 => n18816, B2 => 
                           n23909, ZN => n16339);
   U15367 : OAI22_X1 port map( A1 => n18807, A2 => n23918, B1 => n18871, B2 => 
                           n23909, ZN => n16318);
   U15368 : OAI22_X1 port map( A1 => n18753, A2 => n23918, B1 => n18817, B2 => 
                           n23909, ZN => n16297);
   U15369 : OAI22_X1 port map( A1 => n18806, A2 => n23919, B1 => n18870, B2 => 
                           n23910, ZN => n16276);
   U15370 : OAI22_X1 port map( A1 => n18754, A2 => n23919, B1 => n18818, B2 => 
                           n23910, ZN => n16255);
   U15371 : OAI22_X1 port map( A1 => n18805, A2 => n23919, B1 => n18869, B2 => 
                           n23910, ZN => n16234);
   U15372 : OAI22_X1 port map( A1 => n18755, A2 => n23919, B1 => n18819, B2 => 
                           n23910, ZN => n16213);
   U15373 : OAI22_X1 port map( A1 => n18804, A2 => n23919, B1 => n18868, B2 => 
                           n23910, ZN => n16192);
   U15374 : OAI22_X1 port map( A1 => n18756, A2 => n23919, B1 => n18820, B2 => 
                           n23910, ZN => n16171);
   U15375 : OAI22_X1 port map( A1 => n18803, A2 => n23919, B1 => n18867, B2 => 
                           n23910, ZN => n16150);
   U15376 : OAI22_X1 port map( A1 => n18757, A2 => n23919, B1 => n18821, B2 => 
                           n23910, ZN => n16129);
   U15377 : OAI22_X1 port map( A1 => n18802, A2 => n23919, B1 => n18866, B2 => 
                           n23910, ZN => n16108);
   U15378 : OAI22_X1 port map( A1 => n18758, A2 => n23919, B1 => n18822, B2 => 
                           n23910, ZN => n16087);
   U15379 : OAI22_X1 port map( A1 => n18801, A2 => n23919, B1 => n18865, B2 => 
                           n23910, ZN => n16066);
   U15380 : OAI22_X1 port map( A1 => n18759, A2 => n23919, B1 => n18823, B2 => 
                           n23910, ZN => n16045);
   U15381 : OAI22_X1 port map( A1 => n18800, A2 => n23920, B1 => n18864, B2 => 
                           n23911, ZN => n16024);
   U15382 : OAI22_X1 port map( A1 => n18760, A2 => n23920, B1 => n18824, B2 => 
                           n23911, ZN => n16003);
   U15383 : OAI22_X1 port map( A1 => n18799, A2 => n23920, B1 => n18863, B2 => 
                           n23911, ZN => n15982);
   U15384 : OAI22_X1 port map( A1 => n18761, A2 => n23920, B1 => n18825, B2 => 
                           n23911, ZN => n15961);
   U15385 : OAI22_X1 port map( A1 => n18798, A2 => n23920, B1 => n18862, B2 => 
                           n23911, ZN => n15940);
   U15386 : OAI22_X1 port map( A1 => n18762, A2 => n23920, B1 => n18826, B2 => 
                           n23911, ZN => n15919);
   U15387 : OAI22_X1 port map( A1 => n18797, A2 => n23920, B1 => n18861, B2 => 
                           n23911, ZN => n15898);
   U15388 : OAI22_X1 port map( A1 => n18763, A2 => n23920, B1 => n18827, B2 => 
                           n23911, ZN => n15877);
   U15389 : OAI22_X1 port map( A1 => n18796, A2 => n23920, B1 => n18860, B2 => 
                           n23911, ZN => n15856);
   U15390 : OAI22_X1 port map( A1 => n18764, A2 => n23920, B1 => n18828, B2 => 
                           n23911, ZN => n15835);
   U15391 : OAI22_X1 port map( A1 => n18795, A2 => n23920, B1 => n18859, B2 => 
                           n23911, ZN => n15814);
   U15392 : OAI22_X1 port map( A1 => n18765, A2 => n23920, B1 => n18829, B2 => 
                           n23911, ZN => n15793);
   U15393 : OAI22_X1 port map( A1 => n18794, A2 => n23921, B1 => n18858, B2 => 
                           n23912, ZN => n15772);
   U15394 : OAI22_X1 port map( A1 => n18766, A2 => n23921, B1 => n18830, B2 => 
                           n23912, ZN => n15751);
   U15395 : OAI22_X1 port map( A1 => n18793, A2 => n23921, B1 => n18857, B2 => 
                           n23912, ZN => n15730);
   U15396 : OAI22_X1 port map( A1 => n18767, A2 => n23921, B1 => n18831, B2 => 
                           n23912, ZN => n15709);
   U15397 : OAI22_X1 port map( A1 => n18792, A2 => n23921, B1 => n18856, B2 => 
                           n23912, ZN => n15688);
   U15398 : OAI22_X1 port map( A1 => n18768, A2 => n23921, B1 => n18832, B2 => 
                           n23912, ZN => n15667);
   U15399 : OAI22_X1 port map( A1 => n18791, A2 => n23921, B1 => n18855, B2 => 
                           n23912, ZN => n15646);
   U15400 : OAI22_X1 port map( A1 => n18769, A2 => n23921, B1 => n18833, B2 => 
                           n23912, ZN => n15625);
   U15401 : OAI22_X1 port map( A1 => n18790, A2 => n23921, B1 => n18854, B2 => 
                           n23912, ZN => n15604);
   U15402 : OAI22_X1 port map( A1 => n18770, A2 => n23921, B1 => n18834, B2 => 
                           n23912, ZN => n15583);
   U15403 : OAI22_X1 port map( A1 => n18789, A2 => n23921, B1 => n18853, B2 => 
                           n23912, ZN => n15562);
   U15404 : OAI22_X1 port map( A1 => n18771, A2 => n23921, B1 => n18835, B2 => 
                           n23912, ZN => n15541);
   U15405 : OAI22_X1 port map( A1 => n18788, A2 => n23922, B1 => n18852, B2 => 
                           n23913, ZN => n15520);
   U15406 : OAI22_X1 port map( A1 => n18772, A2 => n23922, B1 => n18836, B2 => 
                           n23913, ZN => n15499);
   U15407 : OAI22_X1 port map( A1 => n18787, A2 => n23922, B1 => n18851, B2 => 
                           n23913, ZN => n15478);
   U15408 : OAI22_X1 port map( A1 => n18773, A2 => n23922, B1 => n18837, B2 => 
                           n23913, ZN => n15457);
   U15409 : OAI22_X1 port map( A1 => n18786, A2 => n23922, B1 => n18850, B2 => 
                           n23913, ZN => n15436);
   U15410 : OAI22_X1 port map( A1 => n18774, A2 => n23922, B1 => n18838, B2 => 
                           n23913, ZN => n15415);
   U15411 : OAI22_X1 port map( A1 => n18785, A2 => n23922, B1 => n18849, B2 => 
                           n23913, ZN => n15394);
   U15412 : OAI22_X1 port map( A1 => n18775, A2 => n23922, B1 => n18839, B2 => 
                           n23913, ZN => n15373);
   U15413 : OAI22_X1 port map( A1 => n18784, A2 => n23922, B1 => n18848, B2 => 
                           n23913, ZN => n15352);
   U15414 : OAI22_X1 port map( A1 => n18776, A2 => n23922, B1 => n18840, B2 => 
                           n23913, ZN => n15331);
   U15415 : OAI22_X1 port map( A1 => n18783, A2 => n23922, B1 => n18847, B2 => 
                           n23913, ZN => n15310);
   U15416 : OAI22_X1 port map( A1 => n18777, A2 => n23922, B1 => n18841, B2 => 
                           n23913, ZN => n15289);
   U15417 : BUF_X1 port map( A => n15180, Z => n23917);
   U15418 : OAI22_X1 port map( A1 => n18782, A2 => n23923, B1 => n18846, B2 => 
                           n23914, ZN => n15268);
   U15419 : OAI22_X1 port map( A1 => n18778, A2 => n23923, B1 => n18842, B2 => 
                           n23914, ZN => n15247);
   U15420 : OAI22_X1 port map( A1 => n18781, A2 => n23923, B1 => n18845, B2 => 
                           n23914, ZN => n15226);
   U15421 : OAI22_X1 port map( A1 => n18779, A2 => n23923, B1 => n18843, B2 => 
                           n23914, ZN => n15179);
   U15422 : OAI22_X1 port map( A1 => n19512, A2 => n23475, B1 => n19640, B2 => 
                           n23460, ZN => n16995);
   U15423 : OAI22_X1 port map( A1 => n19458, A2 => n23474, B1 => n19586, B2 => 
                           n23459, ZN => n17130);
   U15424 : OAI22_X1 port map( A1 => n19457, A2 => n23474, B1 => n19585, B2 => 
                           n23460, ZN => n17076);
   U15425 : OAI22_X1 port map( A1 => n19456, A2 => n23475, B1 => n19584, B2 => 
                           n23464, ZN => n17022);
   U15426 : OAI22_X1 port map( A1 => n19455, A2 => n23475, B1 => n19583, B2 => 
                           n23462, ZN => n16968);
   U15427 : OAI22_X1 port map( A1 => n19511, A2 => n23475, B1 => n19639, B2 => 
                           n23462, ZN => n17049);
   U15428 : OAI22_X1 port map( A1 => n19459, A2 => n23474, B1 => n19587, B2 => 
                           n23464, ZN => n17184);
   U15429 : OAI22_X1 port map( A1 => n19513, A2 => n23475, B1 => n19641, B2 => 
                           n23461, ZN => n16941);
   U15430 : OAI22_X1 port map( A1 => n19508, A2 => n23474, B1 => n19636, B2 => 
                           n23460, ZN => n17211);
   U15431 : OAI22_X1 port map( A1 => n19509, A2 => n23474, B1 => n19637, B2 => 
                           n23459, ZN => n17157);
   U15432 : OAI22_X1 port map( A1 => n19510, A2 => n23474, B1 => n19638, B2 => 
                           n23463, ZN => n17103);
   U15433 : OAI22_X1 port map( A1 => n19454, A2 => n23475, B1 => n19582, B2 => 
                           n23463, ZN => n16914);
   U15434 : AOI221_X1 port map( B1 => n23444, B2 => n21107, C1 => n23428, C2 =>
                           n21536, A => n16996, ZN => n16993);
   U15435 : AOI221_X1 port map( B1 => n23499, B2 => n21180, C1 => n23483, C2 =>
                           n21592, A => n16995, ZN => n16994);
   U15436 : OAI22_X1 port map( A1 => n19576, A2 => n23421, B1 => n19704, B2 => 
                           n23409, ZN => n16996);
   U15437 : AOI221_X1 port map( B1 => n23444, B2 => n21140, C1 => n23428, C2 =>
                           n21569, A => n17131, ZN => n17128);
   U15438 : AOI221_X1 port map( B1 => n23499, B2 => n21198, C1 => n23483, C2 =>
                           n21625, A => n17130, ZN => n17129);
   U15439 : OAI22_X1 port map( A1 => n19522, A2 => n23420, B1 => n19650, B2 => 
                           n23408, ZN => n17131);
   U15440 : AOI221_X1 port map( B1 => n23444, B2 => n21106, C1 => n23428, C2 =>
                           n21535, A => n17077, ZN => n17074);
   U15441 : AOI221_X1 port map( B1 => n23499, B2 => n21179, C1 => n23483, C2 =>
                           n21591, A => n17076, ZN => n17075);
   U15442 : OAI22_X1 port map( A1 => n19521, A2 => n23420, B1 => n19649, B2 => 
                           n23408, ZN => n17077);
   U15443 : AOI221_X1 port map( B1 => n23444, B2 => n21143, C1 => n23428, C2 =>
                           n21572, A => n17023, ZN => n17020);
   U15444 : AOI221_X1 port map( B1 => n23499, B2 => n21201, C1 => n23483, C2 =>
                           n21628, A => n17022, ZN => n17021);
   U15445 : OAI22_X1 port map( A1 => n19520, A2 => n23421, B1 => n19648, B2 => 
                           n23409, ZN => n17023);
   U15446 : AOI221_X1 port map( B1 => n23444, B2 => n21144, C1 => n23428, C2 =>
                           n21573, A => n16969, ZN => n16966);
   U15447 : AOI221_X1 port map( B1 => n23499, B2 => n21173, C1 => n23483, C2 =>
                           n21629, A => n16968, ZN => n16967);
   U15448 : OAI22_X1 port map( A1 => n19519, A2 => n23421, B1 => n19647, B2 => 
                           n23409, ZN => n16969);
   U15449 : AOI221_X1 port map( B1 => n23444, B2 => n21142, C1 => n23428, C2 =>
                           n21571, A => n17050, ZN => n17047);
   U15450 : AOI221_X1 port map( B1 => n23499, B2 => n21200, C1 => n23483, C2 =>
                           n21627, A => n17049, ZN => n17048);
   U15451 : OAI22_X1 port map( A1 => n19575, A2 => n23421, B1 => n19703, B2 => 
                           n23409, ZN => n17050);
   U15452 : AOI221_X1 port map( B1 => n23445, B2 => n21125, C1 => n23429, C2 =>
                           n21554, A => n17185, ZN => n17182);
   U15453 : AOI221_X1 port map( B1 => n23500, B2 => n21192, C1 => n23484, C2 =>
                           n21610, A => n17184, ZN => n17183);
   U15454 : OAI22_X1 port map( A1 => n19523, A2 => n23420, B1 => n19651, B2 => 
                           n23408, ZN => n17185);
   U15455 : AOI221_X1 port map( B1 => n23443, B2 => n21145, C1 => n23427, C2 =>
                           n21574, A => n16942, ZN => n16939);
   U15456 : AOI221_X1 port map( B1 => n23498, B2 => n21202, C1 => n23482, C2 =>
                           n21630, A => n16941, ZN => n16940);
   U15457 : OAI22_X1 port map( A1 => n19577, A2 => n23421, B1 => n19705, B2 => 
                           n23409, ZN => n16942);
   U15458 : AOI221_X1 port map( B1 => n23445, B2 => n21139, C1 => n23429, C2 =>
                           n21568, A => n17212, ZN => n17209);
   U15459 : AOI221_X1 port map( B1 => n23500, B2 => n21172, C1 => n23484, C2 =>
                           n21624, A => n17211, ZN => n17210);
   U15460 : OAI22_X1 port map( A1 => n19572, A2 => n23420, B1 => n19700, B2 => 
                           n23408, ZN => n17212);
   U15461 : AOI221_X1 port map( B1 => n23445, B2 => n21105, C1 => n23429, C2 =>
                           n21534, A => n17158, ZN => n17155);
   U15462 : AOI221_X1 port map( B1 => n23500, B2 => n21178, C1 => n23484, C2 =>
                           n21590, A => n17157, ZN => n17156);
   U15463 : OAI22_X1 port map( A1 => n19573, A2 => n23420, B1 => n19701, B2 => 
                           n23408, ZN => n17158);
   U15464 : AOI221_X1 port map( B1 => n23444, B2 => n21141, C1 => n23428, C2 =>
                           n21570, A => n17104, ZN => n17101);
   U15465 : AOI221_X1 port map( B1 => n23499, B2 => n21199, C1 => n23483, C2 =>
                           n21626, A => n17103, ZN => n17102);
   U15466 : OAI22_X1 port map( A1 => n19574, A2 => n23420, B1 => n19702, B2 => 
                           n23408, ZN => n17104);
   U15467 : AOI221_X1 port map( B1 => n23443, B2 => n21108, C1 => n23427, C2 =>
                           n21537, A => n16915, ZN => n16912);
   U15468 : AOI221_X1 port map( B1 => n23498, B2 => n21181, C1 => n23482, C2 =>
                           n21593, A => n16914, ZN => n16913);
   U15469 : OAI22_X1 port map( A1 => n19518, A2 => n23421, B1 => n19646, B2 => 
                           n23409, ZN => n16915);
   U15470 : OAI22_X1 port map( A1 => n19495, A2 => n23471, B1 => n19623, B2 => 
                           n23461, ZN => n17913);
   U15471 : AOI221_X1 port map( B1 => n23449, B2 => n21208, C1 => n23433, C2 =>
                           n21637, A => n17914, ZN => n17911);
   U15472 : AOI221_X1 port map( B1 => n23504, B2 => n21209, C1 => n23488, C2 =>
                           n21638, A => n17913, ZN => n17912);
   U15473 : OAI22_X1 port map( A1 => n19559, A2 => n23420, B1 => n19687, B2 => 
                           n23406, ZN => n17914);
   U15474 : OAI22_X1 port map( A1 => n19000, A2 => n23475, B1 => n19128, B2 => 
                           n23460, ZN => n16991);
   U15475 : OAI22_X1 port map( A1 => n18946, A2 => n23474, B1 => n19074, B2 => 
                           n23460, ZN => n17126);
   U15476 : OAI22_X1 port map( A1 => n18945, A2 => n23474, B1 => n19073, B2 => 
                           n23461, ZN => n17072);
   U15477 : OAI22_X1 port map( A1 => n18944, A2 => n23475, B1 => n19072, B2 => 
                           n23461, ZN => n17018);
   U15478 : OAI22_X1 port map( A1 => n18943, A2 => n23475, B1 => n19071, B2 => 
                           n23462, ZN => n16964);
   U15479 : OAI22_X1 port map( A1 => n18999, A2 => n23475, B1 => n19127, B2 => 
                           n23463, ZN => n17045);
   U15480 : OAI22_X1 port map( A1 => n18947, A2 => n23474, B1 => n19075, B2 => 
                           n23463, ZN => n17180);
   U15481 : OAI22_X1 port map( A1 => n19001, A2 => n23475, B1 => n19129, B2 => 
                           n23459, ZN => n16937);
   U15482 : OAI22_X1 port map( A1 => n18996, A2 => n23474, B1 => n19124, B2 => 
                           n23461, ZN => n17207);
   U15483 : OAI22_X1 port map( A1 => n18997, A2 => n23474, B1 => n19125, B2 => 
                           n23464, ZN => n17153);
   U15484 : OAI22_X1 port map( A1 => n18998, A2 => n23474, B1 => n19126, B2 => 
                           n23462, ZN => n17099);
   U15485 : OAI22_X1 port map( A1 => n18942, A2 => n23475, B1 => n19070, B2 => 
                           n23459, ZN => n16910);
   U15486 : AOI221_X1 port map( B1 => n23444, B2 => n20912, C1 => n23428, C2 =>
                           n21652, A => n16992, ZN => n16989);
   U15487 : AOI221_X1 port map( B1 => n23499, B2 => n21223, C1 => n23483, C2 =>
                           n21708, A => n16991, ZN => n16990);
   U15488 : OAI22_X1 port map( A1 => n19064, A2 => n23421, B1 => n19192, B2 => 
                           n23409, ZN => n16992);
   U15489 : AOI221_X1 port map( B1 => n23444, B2 => n20946, C1 => n23428, C2 =>
                           n21686, A => n17127, ZN => n17124);
   U15490 : AOI221_X1 port map( B1 => n23499, B2 => n21258, C1 => n23483, C2 =>
                           n21742, A => n17126, ZN => n17125);
   U15491 : OAI22_X1 port map( A1 => n19010, A2 => n23420, B1 => n19138, B2 => 
                           n23408, ZN => n17127);
   U15492 : AOI221_X1 port map( B1 => n23444, B2 => n20911, C1 => n23428, C2 =>
                           n21651, A => n17073, ZN => n17070);
   U15493 : AOI221_X1 port map( B1 => n23499, B2 => n21222, C1 => n23483, C2 =>
                           n21707, A => n17072, ZN => n17071);
   U15494 : OAI22_X1 port map( A1 => n19009, A2 => n23420, B1 => n19137, B2 => 
                           n23408, ZN => n17073);
   U15495 : AOI221_X1 port map( B1 => n23444, B2 => n20949, C1 => n23428, C2 =>
                           n21689, A => n17019, ZN => n17016);
   U15496 : AOI221_X1 port map( B1 => n23499, B2 => n21243, C1 => n23483, C2 =>
                           n21745, A => n17018, ZN => n17017);
   U15497 : OAI22_X1 port map( A1 => n19008, A2 => n23421, B1 => n19136, B2 => 
                           n23409, ZN => n17019);
   U15498 : AOI221_X1 port map( B1 => n23443, B2 => n20950, C1 => n23427, C2 =>
                           n21690, A => n16965, ZN => n16962);
   U15499 : AOI221_X1 port map( B1 => n23498, B2 => n21261, C1 => n23482, C2 =>
                           n21746, A => n16964, ZN => n16963);
   U15500 : OAI22_X1 port map( A1 => n19007, A2 => n23421, B1 => n19135, B2 => 
                           n23409, ZN => n16965);
   U15501 : AOI221_X1 port map( B1 => n23444, B2 => n20948, C1 => n23428, C2 =>
                           n21688, A => n17046, ZN => n17043);
   U15502 : AOI221_X1 port map( B1 => n23499, B2 => n21260, C1 => n23483, C2 =>
                           n21744, A => n17045, ZN => n17044);
   U15503 : OAI22_X1 port map( A1 => n19063, A2 => n23421, B1 => n19191, B2 => 
                           n23409, ZN => n17046);
   U15504 : AOI221_X1 port map( B1 => n23445, B2 => n20930, C1 => n23429, C2 =>
                           n21670, A => n17181, ZN => n17178);
   U15505 : AOI221_X1 port map( B1 => n23500, B2 => n21241, C1 => n23484, C2 =>
                           n21726, A => n17180, ZN => n17179);
   U15506 : OAI22_X1 port map( A1 => n19011, A2 => n23420, B1 => n19139, B2 => 
                           n23408, ZN => n17181);
   U15507 : AOI221_X1 port map( B1 => n23443, B2 => n20951, C1 => n23427, C2 =>
                           n21691, A => n16938, ZN => n16935);
   U15508 : AOI221_X1 port map( B1 => n23498, B2 => n21262, C1 => n23482, C2 =>
                           n21747, A => n16937, ZN => n16936);
   U15509 : OAI22_X1 port map( A1 => n19065, A2 => n23421, B1 => n19193, B2 => 
                           n23409, ZN => n16938);
   U15510 : AOI221_X1 port map( B1 => n23445, B2 => n20945, C1 => n23429, C2 =>
                           n21685, A => n17208, ZN => n17205);
   U15511 : AOI221_X1 port map( B1 => n23500, B2 => n21257, C1 => n23484, C2 =>
                           n21741, A => n17207, ZN => n17206);
   U15512 : OAI22_X1 port map( A1 => n19060, A2 => n23420, B1 => n19188, B2 => 
                           n23408, ZN => n17208);
   U15513 : AOI221_X1 port map( B1 => n23445, B2 => n20910, C1 => n23429, C2 =>
                           n21650, A => n17154, ZN => n17151);
   U15514 : AOI221_X1 port map( B1 => n23500, B2 => n21221, C1 => n23484, C2 =>
                           n21706, A => n17153, ZN => n17152);
   U15515 : OAI22_X1 port map( A1 => n19061, A2 => n23420, B1 => n19189, B2 => 
                           n23408, ZN => n17154);
   U15516 : AOI221_X1 port map( B1 => n23444, B2 => n20947, C1 => n23428, C2 =>
                           n21687, A => n17100, ZN => n17097);
   U15517 : AOI221_X1 port map( B1 => n23499, B2 => n21259, C1 => n23483, C2 =>
                           n21743, A => n17099, ZN => n17098);
   U15518 : OAI22_X1 port map( A1 => n19062, A2 => n23420, B1 => n19190, B2 => 
                           n23408, ZN => n17100);
   U15519 : AOI221_X1 port map( B1 => n23443, B2 => n20913, C1 => n23427, C2 =>
                           n21653, A => n16911, ZN => n16908);
   U15520 : AOI221_X1 port map( B1 => n23498, B2 => n21224, C1 => n23482, C2 =>
                           n21709, A => n16910, ZN => n16909);
   U15521 : OAI22_X1 port map( A1 => n19006, A2 => n23421, B1 => n19134, B2 => 
                           n23409, ZN => n16911);
   U15522 : OAI22_X1 port map( A1 => n19514, A2 => n23471, B1 => n19642, B2 => 
                           n23464, ZN => n16887);
   U15523 : OAI22_X1 port map( A1 => n19453, A2 => n23471, B1 => n19581, B2 => 
                           n23464, ZN => n16860);
   U15524 : OAI22_X1 port map( A1 => n19515, A2 => n23475, B1 => n19643, B2 => 
                           n23464, ZN => n16833);
   U15525 : OAI22_X1 port map( A1 => n19452, A2 => n23472, B1 => n19580, B2 => 
                           n23464, ZN => n16790);
   U15526 : AOI221_X1 port map( B1 => n23443, B2 => n21147, C1 => n23427, C2 =>
                           n21576, A => n16888, ZN => n16885);
   U15527 : AOI221_X1 port map( B1 => n23498, B2 => n21204, C1 => n23482, C2 =>
                           n21633, A => n16887, ZN => n16886);
   U15528 : OAI22_X1 port map( A1 => n19578, A2 => n23417, B1 => n19706, B2 => 
                           n23410, ZN => n16888);
   U15529 : AOI221_X1 port map( B1 => n23443, B2 => n21148, C1 => n23427, C2 =>
                           n21577, A => n16861, ZN => n16858);
   U15530 : AOI221_X1 port map( B1 => n23498, B2 => n21205, C1 => n23482, C2 =>
                           n21634, A => n16860, ZN => n16859);
   U15531 : OAI22_X1 port map( A1 => n19517, A2 => n23419, B1 => n19645, B2 => 
                           n23410, ZN => n16861);
   U15532 : AOI221_X1 port map( B1 => n23443, B2 => n21146, C1 => n23427, C2 =>
                           n21575, A => n16834, ZN => n16831);
   U15533 : AOI221_X1 port map( B1 => n23498, B2 => n21203, C1 => n23482, C2 =>
                           n21632, A => n16833, ZN => n16832);
   U15534 : OAI22_X1 port map( A1 => n19579, A2 => n23416, B1 => n19707, B2 => 
                           n23410, ZN => n16834);
   U15535 : AOI221_X1 port map( B1 => n23443, B2 => n21149, C1 => n23427, C2 =>
                           n21578, A => n16791, ZN => n16787);
   U15536 : AOI221_X1 port map( B1 => n23498, B2 => n21206, C1 => n23482, C2 =>
                           n21635, A => n16790, ZN => n16788);
   U15537 : OAI22_X1 port map( A1 => n19516, A2 => n23416, B1 => n19644, B2 => 
                           n23410, ZN => n16791);
   U15538 : OAI22_X1 port map( A1 => n19466, A2 => n23472, B1 => n19594, B2 => 
                           n23464, ZN => n17562);
   U15539 : OAI22_X1 port map( A1 => n19506, A2 => n23473, B1 => n19634, B2 => 
                           n23463, ZN => n17319);
   U15540 : OAI22_X1 port map( A1 => n19503, A2 => n23473, B1 => n19631, B2 => 
                           n23462, ZN => n17481);
   U15541 : OAI22_X1 port map( A1 => n19460, A2 => n23473, B1 => n19588, B2 => 
                           n23463, ZN => n17238);
   U15542 : OAI22_X1 port map( A1 => n19500, A2 => n23475, B1 => n19628, B2 => 
                           n23460, ZN => n17643);
   U15543 : OAI22_X1 port map( A1 => n19467, A2 => n23473, B1 => n19595, B2 => 
                           n23460, ZN => n17616);
   U15544 : OAI22_X1 port map( A1 => n19464, A2 => n23473, B1 => n19592, B2 => 
                           n23462, ZN => n17454);
   U15545 : OAI22_X1 port map( A1 => n19463, A2 => n23472, B1 => n19591, B2 => 
                           n23462, ZN => n17400);
   U15546 : OAI22_X1 port map( A1 => n19505, A2 => n23473, B1 => n19633, B2 => 
                           n23463, ZN => n17373);
   U15547 : OAI22_X1 port map( A1 => n19461, A2 => n23473, B1 => n19589, B2 => 
                           n23463, ZN => n17292);
   U15548 : OAI22_X1 port map( A1 => n19462, A2 => n23473, B1 => n19590, B2 => 
                           n23463, ZN => n17346);
   U15549 : OAI22_X1 port map( A1 => n19507, A2 => n23473, B1 => n19635, B2 => 
                           n23463, ZN => n17265);
   U15550 : OAI22_X1 port map( A1 => n19502, A2 => n23475, B1 => n19630, B2 => 
                           n23462, ZN => n17535);
   U15551 : OAI22_X1 port map( A1 => n19504, A2 => n23475, B1 => n19632, B2 => 
                           n23462, ZN => n17427);
   U15552 : AOI221_X1 port map( B1 => n23447, B2 => n21100, C1 => n23431, C2 =>
                           n21529, A => n17563, ZN => n17560);
   U15553 : AOI221_X1 port map( B1 => n23502, B2 => n21154, C1 => n23486, C2 =>
                           n21585, A => n17562, ZN => n17561);
   U15554 : OAI22_X1 port map( A1 => n19530, A2 => n23418, B1 => n19658, B2 => 
                           n23410, ZN => n17563);
   U15555 : AOI221_X1 port map( B1 => n23446, B2 => n21103, C1 => n23430, C2 =>
                           n21532, A => n17320, ZN => n17317);
   U15556 : AOI221_X1 port map( B1 => n23501, B2 => n21157, C1 => n23485, C2 =>
                           n21588, A => n17319, ZN => n17318);
   U15557 : OAI22_X1 port map( A1 => n19570, A2 => n23419, B1 => n19698, B2 => 
                           n23409, ZN => n17320);
   U15558 : AOI221_X1 port map( B1 => n23446, B2 => n21124, C1 => n23430, C2 =>
                           n21553, A => n17482, ZN => n17479);
   U15559 : AOI221_X1 port map( B1 => n23501, B2 => n21191, C1 => n23485, C2 =>
                           n21609, A => n17481, ZN => n17480);
   U15560 : OAI22_X1 port map( A1 => n19567, A2 => n23418, B1 => n19695, B2 => 
                           n23407, ZN => n17482);
   U15561 : AOI221_X1 port map( B1 => n23445, B2 => n21104, C1 => n23429, C2 =>
                           n21533, A => n17239, ZN => n17236);
   U15562 : AOI221_X1 port map( B1 => n23500, B2 => n21177, C1 => n23484, C2 =>
                           n21589, A => n17238, ZN => n17237);
   U15563 : OAI22_X1 port map( A1 => n19524, A2 => n23419, B1 => n19652, B2 => 
                           n23408, ZN => n17239);
   U15564 : AOI221_X1 port map( B1 => n23447, B2 => n21269, C1 => n23431, C2 =>
                           n21755, A => n17644, ZN => n17641);
   U15565 : AOI221_X1 port map( B1 => n23502, B2 => n21275, C1 => n23486, C2 =>
                           n21760, A => n17643, ZN => n17642);
   U15566 : OAI22_X1 port map( A1 => n19564, A2 => n23418, B1 => n19692, B2 => 
                           n23405, ZN => n17644);
   U15567 : AOI221_X1 port map( B1 => n23447, B2 => n21099, C1 => n23431, C2 =>
                           n21528, A => n17617, ZN => n17614);
   U15568 : AOI221_X1 port map( B1 => n23502, B2 => n21153, C1 => n23486, C2 =>
                           n21584, A => n17616, ZN => n17615);
   U15569 : OAI22_X1 port map( A1 => n19531, A2 => n23418, B1 => n19659, B2 => 
                           n23405, ZN => n17617);
   U15570 : AOI221_X1 port map( B1 => n23446, B2 => n21101, C1 => n23430, C2 =>
                           n21530, A => n17455, ZN => n17452);
   U15571 : AOI221_X1 port map( B1 => n23501, B2 => n21155, C1 => n23485, C2 =>
                           n21586, A => n17454, ZN => n17453);
   U15572 : OAI22_X1 port map( A1 => n19528, A2 => n23419, B1 => n19656, B2 => 
                           n23406, ZN => n17455);
   U15573 : AOI221_X1 port map( B1 => n23446, B2 => n21135, C1 => n23430, C2 =>
                           n21564, A => n17401, ZN => n17398);
   U15574 : AOI221_X1 port map( B1 => n23501, B2 => n21169, C1 => n23485, C2 =>
                           n21620, A => n17400, ZN => n17399);
   U15575 : OAI22_X1 port map( A1 => n19527, A2 => n23418, B1 => n19655, B2 => 
                           n23405, ZN => n17401);
   U15576 : AOI221_X1 port map( B1 => n23446, B2 => n21102, C1 => n23430, C2 =>
                           n21531, A => n17374, ZN => n17371);
   U15577 : AOI221_X1 port map( B1 => n23501, B2 => n21156, C1 => n23485, C2 =>
                           n21587, A => n17373, ZN => n17372);
   U15578 : OAI22_X1 port map( A1 => n19569, A2 => n23419, B1 => n19697, B2 => 
                           n23409, ZN => n17374);
   U15579 : AOI221_X1 port map( B1 => n23445, B2 => n21137, C1 => n23429, C2 =>
                           n21566, A => n17293, ZN => n17290);
   U15580 : AOI221_X1 port map( B1 => n23500, B2 => n21197, C1 => n23484, C2 =>
                           n21622, A => n17292, ZN => n17291);
   U15581 : OAI22_X1 port map( A1 => n19525, A2 => n23419, B1 => n19653, B2 => 
                           n23406, ZN => n17293);
   U15582 : AOI221_X1 port map( B1 => n23446, B2 => n21136, C1 => n23430, C2 =>
                           n21565, A => n17347, ZN => n17344);
   U15583 : AOI221_X1 port map( B1 => n23501, B2 => n21170, C1 => n23485, C2 =>
                           n21621, A => n17346, ZN => n17345);
   U15584 : OAI22_X1 port map( A1 => n19526, A2 => n23419, B1 => n19654, B2 => 
                           n23405, ZN => n17347);
   U15585 : AOI221_X1 port map( B1 => n23445, B2 => n21138, C1 => n23429, C2 =>
                           n21567, A => n17266, ZN => n17263);
   U15586 : AOI221_X1 port map( B1 => n23500, B2 => n21171, C1 => n23484, C2 =>
                           n21623, A => n17265, ZN => n17264);
   U15587 : OAI22_X1 port map( A1 => n19571, A2 => n23419, B1 => n19699, B2 => 
                           n23407, ZN => n17266);
   U15588 : AOI221_X1 port map( B1 => n23447, B2 => n21270, C1 => n23431, C2 =>
                           n21756, A => n17536, ZN => n17533);
   U15589 : AOI221_X1 port map( B1 => n23502, B2 => n21276, C1 => n23486, C2 =>
                           n21761, A => n17535, ZN => n17534);
   U15590 : OAI22_X1 port map( A1 => n19566, A2 => n23416, B1 => n19694, B2 => 
                           n23410, ZN => n17536);
   U15591 : AOI221_X1 port map( B1 => n23446, B2 => n21268, C1 => n23430, C2 =>
                           n21753, A => n17428, ZN => n17425);
   U15592 : AOI221_X1 port map( B1 => n23501, B2 => n21273, C1 => n23485, C2 =>
                           n21759, A => n17427, ZN => n17426);
   U15593 : OAI22_X1 port map( A1 => n19568, A2 => n23421, B1 => n19696, B2 => 
                           n23407, ZN => n17428);
   U15594 : OAI22_X1 port map( A1 => n19474, A2 => n23473, B1 => n19602, B2 => 
                           n23461, ZN => n17994);
   U15595 : OAI22_X1 port map( A1 => n19499, A2 => n23471, B1 => n19627, B2 => 
                           n23459, ZN => n17697);
   U15596 : OAI22_X1 port map( A1 => n19472, A2 => n23474, B1 => n19600, B2 => 
                           n23461, ZN => n17886);
   U15597 : OAI22_X1 port map( A1 => n19469, A2 => n23472, B1 => n19597, B2 => 
                           n23462, ZN => n17724);
   U15598 : OAI22_X1 port map( A1 => n19468, A2 => n23475, B1 => n19596, B2 => 
                           n23463, ZN => n17670);
   U15599 : OAI22_X1 port map( A1 => n19497, A2 => n23472, B1 => n19625, B2 => 
                           n23461, ZN => n17805);
   U15600 : OAI22_X1 port map( A1 => n19498, A2 => n23472, B1 => n19626, B2 => 
                           n23464, ZN => n17751);
   U15601 : OAI22_X1 port map( A1 => n19493, A2 => n23475, B1 => n19621, B2 => 
                           n23461, ZN => n18021);
   U15602 : OAI22_X1 port map( A1 => n19501, A2 => n23473, B1 => n19629, B2 => 
                           n23462, ZN => n17589);
   U15603 : OAI22_X1 port map( A1 => n19494, A2 => n23472, B1 => n19622, B2 => 
                           n23461, ZN => n17967);
   U15604 : OAI22_X1 port map( A1 => n19470, A2 => n23472, B1 => n19598, B2 => 
                           n23463, ZN => n17778);
   U15605 : OAI22_X1 port map( A1 => n19496, A2 => n23472, B1 => n19624, B2 => 
                           n23464, ZN => n17859);
   U15606 : OAI22_X1 port map( A1 => n19473, A2 => n23474, B1 => n19601, B2 => 
                           n23461, ZN => n17940);
   U15607 : OAI22_X1 port map( A1 => n19471, A2 => n23472, B1 => n19599, B2 => 
                           n23459, ZN => n17832);
   U15608 : AOI221_X1 port map( B1 => n23449, B2 => n21096, C1 => n23433, C2 =>
                           n21525, A => n17995, ZN => n17992);
   U15609 : AOI221_X1 port map( B1 => n23504, B2 => n21152, C1 => n23488, C2 =>
                           n21581, A => n17994, ZN => n17993);
   U15610 : OAI22_X1 port map( A1 => n19538, A2 => n23419, B1 => n19666, B2 => 
                           n23406, ZN => n17995);
   U15611 : AOI221_X1 port map( B1 => n23448, B2 => n21122, C1 => n23432, C2 =>
                           n21551, A => n17698, ZN => n17695);
   U15612 : AOI221_X1 port map( B1 => n23503, B2 => n21190, C1 => n23487, C2 =>
                           n21607, A => n17697, ZN => n17696);
   U15613 : OAI22_X1 port map( A1 => n19563, A2 => n23418, B1 => n19691, B2 => 
                           n23410, ZN => n17698);
   U15614 : AOI221_X1 port map( B1 => n23449, B2 => n21119, C1 => n23433, C2 =>
                           n21548, A => n17887, ZN => n17884);
   U15615 : AOI221_X1 port map( B1 => n23504, B2 => n21161, C1 => n23488, C2 =>
                           n21604, A => n17886, ZN => n17885);
   U15616 : OAI22_X1 port map( A1 => n19536, A2 => n23418, B1 => n19664, B2 => 
                           n23406, ZN => n17887);
   U15617 : AOI221_X1 port map( B1 => n23448, B2 => n21121, C1 => n23432, C2 =>
                           n21550, A => n17725, ZN => n17722);
   U15618 : AOI221_X1 port map( B1 => n23503, B2 => n21189, C1 => n23487, C2 =>
                           n21606, A => n17724, ZN => n17723);
   U15619 : OAI22_X1 port map( A1 => n19533, A2 => n23417, B1 => n19661, B2 => 
                           n23407, ZN => n17725);
   U15620 : AOI221_X1 port map( B1 => n23448, B2 => n21123, C1 => n23432, C2 =>
                           n21552, A => n17671, ZN => n17668);
   U15621 : AOI221_X1 port map( B1 => n23503, B2 => n21163, C1 => n23487, C2 =>
                           n21608, A => n17670, ZN => n17669);
   U15622 : OAI22_X1 port map( A1 => n19532, A2 => n23418, B1 => n19660, B2 => 
                           n23408, ZN => n17671);
   U15623 : AOI221_X1 port map( B1 => n23448, B2 => n21098, C1 => n23432, C2 =>
                           n21527, A => n17806, ZN => n17803);
   U15624 : AOI221_X1 port map( B1 => n23503, B2 => n21176, C1 => n23487, C2 =>
                           n21583, A => n17805, ZN => n17804);
   U15625 : OAI22_X1 port map( A1 => n19561, A2 => n23417, B1 => n19689, B2 => 
                           n23407, ZN => n17806);
   U15626 : AOI221_X1 port map( B1 => n23448, B2 => n21133, C1 => n23432, C2 =>
                           n21562, A => n17752, ZN => n17749);
   U15627 : AOI221_X1 port map( B1 => n23503, B2 => n21196, C1 => n23487, C2 =>
                           n21618, A => n17751, ZN => n17750);
   U15628 : OAI22_X1 port map( A1 => n19562, A2 => n23417, B1 => n19690, B2 => 
                           n23407, ZN => n17752);
   U15629 : AOI221_X1 port map( B1 => n23450, B2 => n21117, C1 => n23434, C2 =>
                           n21546, A => n18022, ZN => n18019);
   U15630 : AOI221_X1 port map( B1 => n23505, B2 => n21160, C1 => n23489, C2 =>
                           n21602, A => n18021, ZN => n18020);
   U15631 : OAI22_X1 port map( A1 => n19557, A2 => n23421, B1 => n19685, B2 => 
                           n23406, ZN => n18022);
   U15632 : AOI221_X1 port map( B1 => n23447, B2 => n21134, C1 => n23431, C2 =>
                           n21563, A => n17590, ZN => n17587);
   U15633 : AOI221_X1 port map( B1 => n23502, B2 => n21168, C1 => n23486, C2 =>
                           n21619, A => n17589, ZN => n17588);
   U15634 : OAI22_X1 port map( A1 => n19565, A2 => n23418, B1 => n19693, B2 => 
                           n23409, ZN => n17590);
   U15635 : AOI221_X1 port map( B1 => n23449, B2 => n21118, C1 => n23433, C2 =>
                           n21547, A => n17968, ZN => n17965);
   U15636 : AOI221_X1 port map( B1 => n23504, B2 => n21188, C1 => n23488, C2 =>
                           n21603, A => n17967, ZN => n17966);
   U15637 : OAI22_X1 port map( A1 => n19558, A2 => n23417, B1 => n19686, B2 => 
                           n23406, ZN => n17968);
   U15638 : AOI221_X1 port map( B1 => n23448, B2 => n21120, C1 => n23432, C2 =>
                           n21549, A => n17779, ZN => n17776);
   U15639 : AOI221_X1 port map( B1 => n23503, B2 => n21162, C1 => n23487, C2 =>
                           n21605, A => n17778, ZN => n17777);
   U15640 : OAI22_X1 port map( A1 => n19534, A2 => n23417, B1 => n19662, B2 => 
                           n23407, ZN => n17779);
   U15641 : AOI221_X1 port map( B1 => n23449, B2 => n21097, C1 => n23433, C2 =>
                           n21526, A => n17860, ZN => n17857);
   U15642 : AOI221_X1 port map( B1 => n23504, B2 => n21175, C1 => n23488, C2 =>
                           n21582, A => n17859, ZN => n17858);
   U15643 : OAI22_X1 port map( A1 => n19560, A2 => n23417, B1 => n19688, B2 => 
                           n23407, ZN => n17860);
   U15644 : AOI221_X1 port map( B1 => n23449, B2 => n21131, C1 => n23433, C2 =>
                           n21560, A => n17941, ZN => n17938);
   U15645 : AOI221_X1 port map( B1 => n23504, B2 => n21167, C1 => n23488, C2 =>
                           n21616, A => n17940, ZN => n17939);
   U15646 : OAI22_X1 port map( A1 => n19537, A2 => n23420, B1 => n19665, B2 => 
                           n23406, ZN => n17941);
   U15647 : AOI221_X1 port map( B1 => n23449, B2 => n21132, C1 => n23433, C2 =>
                           n21561, A => n17833, ZN => n17830);
   U15648 : AOI221_X1 port map( B1 => n23504, B2 => n21195, C1 => n23488, C2 =>
                           n21617, A => n17832, ZN => n17831);
   U15649 : OAI22_X1 port map( A1 => n19535, A2 => n23417, B1 => n19663, B2 => 
                           n23407, ZN => n17833);
   U15650 : OAI22_X1 port map( A1 => n18983, A2 => n23474, B1 => n19111, B2 => 
                           n23461, ZN => n17909);
   U15651 : AOI221_X1 port map( B1 => n23449, B2 => n20956, C1 => n23433, C2 =>
                           n21764, A => n17910, ZN => n17907);
   U15652 : AOI221_X1 port map( B1 => n23504, B2 => n21274, C1 => n23488, C2 =>
                           n21765, A => n17909, ZN => n17908);
   U15653 : OAI22_X1 port map( A1 => n19047, A2 => n23416, B1 => n19175, B2 => 
                           n23406, ZN => n17910);
   U15654 : OAI22_X1 port map( A1 => n19465, A2 => n23474, B1 => n19593, B2 => 
                           n23462, ZN => n17508);
   U15655 : AOI221_X1 port map( B1 => n23447, B2 => n21271, C1 => n23431, C2 =>
                           n21757, A => n17509, ZN => n17506);
   U15656 : AOI221_X1 port map( B1 => n23502, B2 => n21277, C1 => n23486, C2 =>
                           n21762, A => n17508, ZN => n17507);
   U15657 : OAI22_X1 port map( A1 => n19529, A2 => n23420, B1 => n19657, B2 => 
                           n23410, ZN => n17509);
   U15658 : OAI22_X1 port map( A1 => n19002, A2 => n23472, B1 => n19130, B2 => 
                           n23464, ZN => n16883);
   U15659 : OAI22_X1 port map( A1 => n18941, A2 => n23473, B1 => n19069, B2 => 
                           n23464, ZN => n16856);
   U15660 : OAI22_X1 port map( A1 => n19003, A2 => n23472, B1 => n19131, B2 => 
                           n23464, ZN => n16829);
   U15661 : OAI22_X1 port map( A1 => n18940, A2 => n23471, B1 => n19068, B2 => 
                           n23464, ZN => n16779);
   U15662 : AOI221_X1 port map( B1 => n23443, B2 => n20952, C1 => n23427, C2 =>
                           n21692, A => n16884, ZN => n16881);
   U15663 : AOI221_X1 port map( B1 => n23498, B2 => n21263, C1 => n23482, C2 =>
                           n21748, A => n16883, ZN => n16882);
   U15664 : OAI22_X1 port map( A1 => n19066, A2 => n23416, B1 => n19194, B2 => 
                           n23410, ZN => n16884);
   U15665 : AOI221_X1 port map( B1 => n23443, B2 => n20953, C1 => n23427, C2 =>
                           n21693, A => n16857, ZN => n16854);
   U15666 : AOI221_X1 port map( B1 => n23498, B2 => n21264, C1 => n23482, C2 =>
                           n21749, A => n16856, ZN => n16855);
   U15667 : OAI22_X1 port map( A1 => n19005, A2 => n23421, B1 => n19133, B2 => 
                           n23410, ZN => n16857);
   U15668 : AOI221_X1 port map( B1 => n23443, B2 => n20931, C1 => n23427, C2 =>
                           n21671, A => n16830, ZN => n16827);
   U15669 : AOI221_X1 port map( B1 => n23498, B2 => n21242, C1 => n23482, C2 =>
                           n21727, A => n16829, ZN => n16828);
   U15670 : OAI22_X1 port map( A1 => n19067, A2 => n23417, B1 => n19195, B2 => 
                           n23410, ZN => n16830);
   U15671 : AOI221_X1 port map( B1 => n23448, B2 => n20954, C1 => n23432, C2 =>
                           n21694, A => n16784, ZN => n16774);
   U15672 : AOI221_X1 port map( B1 => n23503, B2 => n21265, C1 => n23487, C2 =>
                           n21750, A => n16779, ZN => n16775);
   U15673 : OAI22_X1 port map( A1 => n19004, A2 => n23419, B1 => n19132, B2 => 
                           n23410, ZN => n16784);
   U15674 : OAI22_X1 port map( A1 => n18954, A2 => n23473, B1 => n19082, B2 => 
                           n23460, ZN => n17558);
   U15675 : OAI22_X1 port map( A1 => n18994, A2 => n23473, B1 => n19122, B2 => 
                           n23463, ZN => n17315);
   U15676 : OAI22_X1 port map( A1 => n18991, A2 => n23475, B1 => n19119, B2 => 
                           n23462, ZN => n17477);
   U15677 : OAI22_X1 port map( A1 => n18948, A2 => n23473, B1 => n19076, B2 => 
                           n23463, ZN => n17234);
   U15678 : OAI22_X1 port map( A1 => n18988, A2 => n23474, B1 => n19116, B2 => 
                           n23459, ZN => n17639);
   U15679 : OAI22_X1 port map( A1 => n18955, A2 => n23471, B1 => n19083, B2 => 
                           n23461, ZN => n17612);
   U15680 : OAI22_X1 port map( A1 => n18952, A2 => n23472, B1 => n19080, B2 => 
                           n23462, ZN => n17450);
   U15681 : OAI22_X1 port map( A1 => n18951, A2 => n23473, B1 => n19079, B2 => 
                           n23462, ZN => n17396);
   U15682 : OAI22_X1 port map( A1 => n18993, A2 => n23473, B1 => n19121, B2 => 
                           n23463, ZN => n17369);
   U15683 : OAI22_X1 port map( A1 => n18949, A2 => n23473, B1 => n19077, B2 => 
                           n23463, ZN => n17288);
   U15684 : OAI22_X1 port map( A1 => n18950, A2 => n23473, B1 => n19078, B2 => 
                           n23463, ZN => n17342);
   U15685 : OAI22_X1 port map( A1 => n18995, A2 => n23473, B1 => n19123, B2 => 
                           n23463, ZN => n17261);
   U15686 : OAI22_X1 port map( A1 => n18990, A2 => n23472, B1 => n19118, B2 => 
                           n23462, ZN => n17531);
   U15687 : OAI22_X1 port map( A1 => n18992, A2 => n23471, B1 => n19120, B2 => 
                           n23462, ZN => n17423);
   U15688 : AOI221_X1 port map( B1 => n23447, B2 => n20905, C1 => n23431, C2 =>
                           n21645, A => n17559, ZN => n17556);
   U15689 : AOI221_X1 port map( B1 => n23502, B2 => n21216, C1 => n23486, C2 =>
                           n21701, A => n17558, ZN => n17557);
   U15690 : OAI22_X1 port map( A1 => n19018, A2 => n23418, B1 => n19146, B2 => 
                           n23409, ZN => n17559);
   U15691 : AOI221_X1 port map( B1 => n23445, B2 => n20908, C1 => n23429, C2 =>
                           n21648, A => n17316, ZN => n17313);
   U15692 : AOI221_X1 port map( B1 => n23500, B2 => n21219, C1 => n23484, C2 =>
                           n21704, A => n17315, ZN => n17314);
   U15693 : OAI22_X1 port map( A1 => n19058, A2 => n23419, B1 => n19186, B2 => 
                           n23410, ZN => n17316);
   U15694 : AOI221_X1 port map( B1 => n23446, B2 => n20929, C1 => n23430, C2 =>
                           n21669, A => n17478, ZN => n17475);
   U15695 : AOI221_X1 port map( B1 => n23501, B2 => n21240, C1 => n23485, C2 =>
                           n21725, A => n17477, ZN => n17476);
   U15696 : OAI22_X1 port map( A1 => n19055, A2 => n23418, B1 => n19183, B2 => 
                           n23405, ZN => n17478);
   U15697 : AOI221_X1 port map( B1 => n23445, B2 => n20909, C1 => n23429, C2 =>
                           n21649, A => n17235, ZN => n17232);
   U15698 : AOI221_X1 port map( B1 => n23500, B2 => n21220, C1 => n23484, C2 =>
                           n21705, A => n17234, ZN => n17233);
   U15699 : OAI22_X1 port map( A1 => n19012, A2 => n23419, B1 => n19140, B2 => 
                           n23407, ZN => n17235);
   U15700 : AOI221_X1 port map( B1 => n23447, B2 => n20959, C1 => n23431, C2 =>
                           n21832, A => n17640, ZN => n17637);
   U15701 : AOI221_X1 port map( B1 => n23502, B2 => n21281, C1 => n23486, C2 =>
                           n21837, A => n17639, ZN => n17638);
   U15702 : OAI22_X1 port map( A1 => n19052, A2 => n23418, B1 => n19180, B2 => 
                           n23405, ZN => n17640);
   U15703 : AOI221_X1 port map( B1 => n23447, B2 => n20904, C1 => n23431, C2 =>
                           n21644, A => n17613, ZN => n17610);
   U15704 : AOI221_X1 port map( B1 => n23502, B2 => n21215, C1 => n23486, C2 =>
                           n21700, A => n17612, ZN => n17611);
   U15705 : OAI22_X1 port map( A1 => n19019, A2 => n23418, B1 => n19147, B2 => 
                           n23408, ZN => n17613);
   U15706 : AOI221_X1 port map( B1 => n23446, B2 => n20906, C1 => n23430, C2 =>
                           n21646, A => n17451, ZN => n17448);
   U15707 : AOI221_X1 port map( B1 => n23501, B2 => n21217, C1 => n23485, C2 =>
                           n21702, A => n17450, ZN => n17449);
   U15708 : OAI22_X1 port map( A1 => n19016, A2 => n23417, B1 => n19144, B2 => 
                           n23407, ZN => n17451);
   U15709 : AOI221_X1 port map( B1 => n23446, B2 => n20941, C1 => n23430, C2 =>
                           n21681, A => n17397, ZN => n17394);
   U15710 : AOI221_X1 port map( B1 => n23501, B2 => n21253, C1 => n23485, C2 =>
                           n21737, A => n17396, ZN => n17395);
   U15711 : OAI22_X1 port map( A1 => n19015, A2 => n23419, B1 => n19143, B2 => 
                           n23408, ZN => n17397);
   U15712 : AOI221_X1 port map( B1 => n23446, B2 => n20907, C1 => n23430, C2 =>
                           n21647, A => n17370, ZN => n17367);
   U15713 : AOI221_X1 port map( B1 => n23501, B2 => n21218, C1 => n23485, C2 =>
                           n21703, A => n17369, ZN => n17368);
   U15714 : OAI22_X1 port map( A1 => n19057, A2 => n23419, B1 => n19185, B2 => 
                           n23406, ZN => n17370);
   U15715 : AOI221_X1 port map( B1 => n23445, B2 => n20943, C1 => n23429, C2 =>
                           n21683, A => n17289, ZN => n17286);
   U15716 : AOI221_X1 port map( B1 => n23500, B2 => n21255, C1 => n23484, C2 =>
                           n21739, A => n17288, ZN => n17287);
   U15717 : OAI22_X1 port map( A1 => n19013, A2 => n23419, B1 => n19141, B2 => 
                           n23407, ZN => n17289);
   U15718 : AOI221_X1 port map( B1 => n23446, B2 => n20942, C1 => n23430, C2 =>
                           n21682, A => n17343, ZN => n17340);
   U15719 : AOI221_X1 port map( B1 => n23501, B2 => n21254, C1 => n23485, C2 =>
                           n21738, A => n17342, ZN => n17341);
   U15720 : OAI22_X1 port map( A1 => n19014, A2 => n23419, B1 => n19142, B2 => 
                           n23409, ZN => n17343);
   U15721 : AOI221_X1 port map( B1 => n23445, B2 => n20944, C1 => n23429, C2 =>
                           n21684, A => n17262, ZN => n17259);
   U15722 : AOI221_X1 port map( B1 => n23500, B2 => n21256, C1 => n23484, C2 =>
                           n21740, A => n17261, ZN => n17260);
   U15723 : OAI22_X1 port map( A1 => n19059, A2 => n23419, B1 => n19187, B2 => 
                           n23410, ZN => n17262);
   U15724 : AOI221_X1 port map( B1 => n23447, B2 => n20960, C1 => n23431, C2 =>
                           n21833, A => n17532, ZN => n17529);
   U15725 : AOI221_X1 port map( B1 => n23502, B2 => n21282, C1 => n23486, C2 =>
                           n21838, A => n17531, ZN => n17530);
   U15726 : OAI22_X1 port map( A1 => n19054, A2 => n23417, B1 => n19182, B2 => 
                           n23405, ZN => n17532);
   U15727 : AOI221_X1 port map( B1 => n23446, B2 => n20958, C1 => n23430, C2 =>
                           n21831, A => n17424, ZN => n17421);
   U15728 : AOI221_X1 port map( B1 => n23501, B2 => n21280, C1 => n23485, C2 =>
                           n21836, A => n17423, ZN => n17422);
   U15729 : OAI22_X1 port map( A1 => n19056, A2 => n23416, B1 => n19184, B2 => 
                           n23406, ZN => n17424);
   U15730 : OAI22_X1 port map( A1 => n18962, A2 => n23472, B1 => n19090, B2 => 
                           n23461, ZN => n17990);
   U15731 : OAI22_X1 port map( A1 => n18987, A2 => n23472, B1 => n19115, B2 => 
                           n23461, ZN => n17693);
   U15732 : OAI22_X1 port map( A1 => n18960, A2 => n23473, B1 => n19088, B2 => 
                           n23461, ZN => n17882);
   U15733 : OAI22_X1 port map( A1 => n18957, A2 => n23472, B1 => n19085, B2 => 
                           n23464, ZN => n17720);
   U15734 : OAI22_X1 port map( A1 => n18956, A2 => n23474, B1 => n19084, B2 => 
                           n23459, ZN => n17666);
   U15735 : OAI22_X1 port map( A1 => n18985, A2 => n23472, B1 => n19113, B2 => 
                           n23462, ZN => n17801);
   U15736 : OAI22_X1 port map( A1 => n18986, A2 => n23472, B1 => n19114, B2 => 
                           n23463, ZN => n17747);
   U15737 : OAI22_X1 port map( A1 => n18981, A2 => n23474, B1 => n19109, B2 => 
                           n23461, ZN => n18017);
   U15738 : OAI22_X1 port map( A1 => n18989, A2 => n23473, B1 => n19117, B2 => 
                           n23464, ZN => n17585);
   U15739 : OAI22_X1 port map( A1 => n18982, A2 => n23472, B1 => n19110, B2 => 
                           n23461, ZN => n17963);
   U15740 : OAI22_X1 port map( A1 => n18958, A2 => n23472, B1 => n19086, B2 => 
                           n23461, ZN => n17774);
   U15741 : OAI22_X1 port map( A1 => n18984, A2 => n23472, B1 => n19112, B2 => 
                           n23463, ZN => n17855);
   U15742 : OAI22_X1 port map( A1 => n18961, A2 => n23475, B1 => n19089, B2 => 
                           n23461, ZN => n17936);
   U15743 : OAI22_X1 port map( A1 => n18959, A2 => n23472, B1 => n19087, B2 => 
                           n23462, ZN => n17828);
   U15744 : AOI221_X1 port map( B1 => n23449, B2 => n20902, C1 => n23433, C2 =>
                           n21642, A => n17991, ZN => n17988);
   U15745 : AOI221_X1 port map( B1 => n23504, B2 => n21212, C1 => n23488, C2 =>
                           n21697, A => n17990, ZN => n17989);
   U15746 : OAI22_X1 port map( A1 => n19026, A2 => n23418, B1 => n19154, B2 => 
                           n23406, ZN => n17991);
   U15747 : AOI221_X1 port map( B1 => n23448, B2 => n20927, C1 => n23432, C2 =>
                           n21667, A => n17694, ZN => n17691);
   U15748 : AOI221_X1 port map( B1 => n23503, B2 => n21238, C1 => n23487, C2 =>
                           n21723, A => n17693, ZN => n17692);
   U15749 : OAI22_X1 port map( A1 => n19051, A2 => n23418, B1 => n19179, B2 => 
                           n23406, ZN => n17694);
   U15750 : AOI221_X1 port map( B1 => n23449, B2 => n20924, C1 => n23433, C2 =>
                           n21664, A => n17883, ZN => n17880);
   U15751 : AOI221_X1 port map( B1 => n23504, B2 => n21235, C1 => n23488, C2 =>
                           n21720, A => n17882, ZN => n17881);
   U15752 : OAI22_X1 port map( A1 => n19024, A2 => n23419, B1 => n19152, B2 => 
                           n23406, ZN => n17883);
   U15753 : AOI221_X1 port map( B1 => n23448, B2 => n20926, C1 => n23432, C2 =>
                           n21666, A => n17721, ZN => n17718);
   U15754 : AOI221_X1 port map( B1 => n23503, B2 => n21237, C1 => n23487, C2 =>
                           n21722, A => n17720, ZN => n17719);
   U15755 : OAI22_X1 port map( A1 => n19021, A2 => n23417, B1 => n19149, B2 => 
                           n23407, ZN => n17721);
   U15756 : AOI221_X1 port map( B1 => n23447, B2 => n20928, C1 => n23431, C2 =>
                           n21668, A => n17667, ZN => n17664);
   U15757 : AOI221_X1 port map( B1 => n23502, B2 => n21239, C1 => n23486, C2 =>
                           n21724, A => n17666, ZN => n17665);
   U15758 : OAI22_X1 port map( A1 => n19020, A2 => n23418, B1 => n19148, B2 => 
                           n23407, ZN => n17667);
   U15759 : AOI221_X1 port map( B1 => n23448, B2 => n20903, C1 => n23432, C2 =>
                           n21643, A => n17802, ZN => n17799);
   U15760 : AOI221_X1 port map( B1 => n23503, B2 => n21214, C1 => n23487, C2 =>
                           n21699, A => n17801, ZN => n17800);
   U15761 : OAI22_X1 port map( A1 => n19049, A2 => n23417, B1 => n19177, B2 => 
                           n23407, ZN => n17802);
   U15762 : AOI221_X1 port map( B1 => n23448, B2 => n20939, C1 => n23432, C2 =>
                           n21679, A => n17748, ZN => n17745);
   U15763 : AOI221_X1 port map( B1 => n23503, B2 => n21251, C1 => n23487, C2 =>
                           n21735, A => n17747, ZN => n17746);
   U15764 : OAI22_X1 port map( A1 => n19050, A2 => n23417, B1 => n19178, B2 => 
                           n23407, ZN => n17748);
   U15765 : AOI221_X1 port map( B1 => n23450, B2 => n20922, C1 => n23434, C2 =>
                           n21662, A => n18018, ZN => n18015);
   U15766 : AOI221_X1 port map( B1 => n23505, B2 => n21233, C1 => n23489, C2 =>
                           n21718, A => n18017, ZN => n18016);
   U15767 : OAI22_X1 port map( A1 => n19045, A2 => n23420, B1 => n19173, B2 => 
                           n23406, ZN => n18018);
   U15768 : AOI221_X1 port map( B1 => n23447, B2 => n20940, C1 => n23431, C2 =>
                           n21680, A => n17586, ZN => n17583);
   U15769 : AOI221_X1 port map( B1 => n23502, B2 => n21252, C1 => n23486, C2 =>
                           n21736, A => n17585, ZN => n17584);
   U15770 : OAI22_X1 port map( A1 => n19053, A2 => n23418, B1 => n19181, B2 => 
                           n23410, ZN => n17586);
   U15771 : AOI221_X1 port map( B1 => n23449, B2 => n20923, C1 => n23433, C2 =>
                           n21663, A => n17964, ZN => n17961);
   U15772 : AOI221_X1 port map( B1 => n23504, B2 => n21234, C1 => n23488, C2 =>
                           n21719, A => n17963, ZN => n17962);
   U15773 : OAI22_X1 port map( A1 => n19046, A2 => n23417, B1 => n19174, B2 => 
                           n23406, ZN => n17964);
   U15774 : AOI221_X1 port map( B1 => n23448, B2 => n20925, C1 => n23432, C2 =>
                           n21665, A => n17775, ZN => n17772);
   U15775 : AOI221_X1 port map( B1 => n23503, B2 => n21236, C1 => n23487, C2 =>
                           n21721, A => n17774, ZN => n17773);
   U15776 : OAI22_X1 port map( A1 => n19022, A2 => n23417, B1 => n19150, B2 => 
                           n23407, ZN => n17775);
   U15777 : AOI221_X1 port map( B1 => n23449, B2 => n20899, C1 => n23433, C2 =>
                           n21639, A => n17856, ZN => n17853);
   U15778 : AOI221_X1 port map( B1 => n23504, B2 => n21213, C1 => n23488, C2 =>
                           n21698, A => n17855, ZN => n17854);
   U15779 : OAI22_X1 port map( A1 => n19048, A2 => n23417, B1 => n19176, B2 => 
                           n23407, ZN => n17856);
   U15780 : AOI221_X1 port map( B1 => n23449, B2 => n20937, C1 => n23433, C2 =>
                           n21677, A => n17937, ZN => n17934);
   U15781 : AOI221_X1 port map( B1 => n23504, B2 => n21249, C1 => n23488, C2 =>
                           n21733, A => n17936, ZN => n17935);
   U15782 : OAI22_X1 port map( A1 => n19025, A2 => n23421, B1 => n19153, B2 => 
                           n23406, ZN => n17937);
   U15783 : AOI221_X1 port map( B1 => n23448, B2 => n20938, C1 => n23432, C2 =>
                           n21678, A => n17829, ZN => n17826);
   U15784 : AOI221_X1 port map( B1 => n23503, B2 => n21250, C1 => n23487, C2 =>
                           n21734, A => n17828, ZN => n17827);
   U15785 : OAI22_X1 port map( A1 => n19023, A2 => n23417, B1 => n19151, B2 => 
                           n23407, ZN => n17829);
   U15786 : OAI22_X1 port map( A1 => n18953, A2 => n23471, B1 => n19081, B2 => 
                           n23462, ZN => n17504);
   U15787 : AOI221_X1 port map( B1 => n23447, B2 => n20961, C1 => n23431, C2 =>
                           n21834, A => n17505, ZN => n17502);
   U15788 : AOI221_X1 port map( B1 => n23502, B2 => n21283, C1 => n23486, C2 =>
                           n21839, A => n17504, ZN => n17503);
   U15789 : OAI22_X1 port map( A1 => n19017, A2 => n23420, B1 => n19145, B2 => 
                           n23409, ZN => n17505);
   U15790 : OAI22_X1 port map( A1 => n19483, A2 => n23471, B1 => n19611, B2 => 
                           n23459, ZN => n18480);
   U15791 : OAI22_X1 port map( A1 => n19482, A2 => n23471, B1 => n19610, B2 => 
                           n23459, ZN => n18426);
   U15792 : OAI22_X1 port map( A1 => n19489, A2 => n23472, B1 => n19617, B2 => 
                           n23460, ZN => n18237);
   U15793 : OAI22_X1 port map( A1 => n19490, A2 => n23471, B1 => n19618, B2 => 
                           n23464, ZN => n18183);
   U15794 : OAI22_X1 port map( A1 => n19486, A2 => n23471, B1 => n19614, B2 => 
                           n23459, ZN => n18399);
   U15795 : OAI22_X1 port map( A1 => n19487, A2 => n23472, B1 => n19615, B2 => 
                           n23460, ZN => n18345);
   U15796 : OAI22_X1 port map( A1 => n19481, A2 => n23471, B1 => n19609, B2 => 
                           n23459, ZN => n18372);
   U15797 : OAI22_X1 port map( A1 => n19478, A2 => n23473, B1 => n19606, B2 => 
                           n23460, ZN => n18210);
   U15798 : OAI22_X1 port map( A1 => n19480, A2 => n23475, B1 => n19608, B2 => 
                           n23460, ZN => n18318);
   U15799 : OAI22_X1 port map( A1 => n19485, A2 => n23471, B1 => n19613, B2 => 
                           n23459, ZN => n18453);
   U15800 : OAI22_X1 port map( A1 => n19479, A2 => n23474, B1 => n19607, B2 => 
                           n23460, ZN => n18264);
   U15801 : OAI22_X1 port map( A1 => n19488, A2 => n23474, B1 => n19616, B2 => 
                           n23460, ZN => n18291);
   U15802 : AOI221_X1 port map( B1 => n23452, B2 => n21094, C1 => n23436, C2 =>
                           n21523, A => n18481, ZN => n18478);
   U15803 : AOI221_X1 port map( B1 => n23507, B2 => n21151, C1 => n23491, C2 =>
                           n21579, A => n18480, ZN => n18479);
   U15804 : OAI22_X1 port map( A1 => n19547, A2 => n23416, B1 => n19675, B2 => 
                           n23405, ZN => n18481);
   U15805 : AOI221_X1 port map( B1 => n23452, B2 => n21110, C1 => n23436, C2 =>
                           n21539, A => n18427, ZN => n18424);
   U15806 : AOI221_X1 port map( B1 => n23507, B2 => n21158, C1 => n23491, C2 =>
                           n21595, A => n18426, ZN => n18425);
   U15807 : OAI22_X1 port map( A1 => n19546, A2 => n23420, B1 => n19674, B2 => 
                           n23409, ZN => n18427);
   U15808 : AOI221_X1 port map( B1 => n23451, B2 => n21128, C1 => n23435, C2 =>
                           n21557, A => n18238, ZN => n18235);
   U15809 : AOI221_X1 port map( B1 => n23506, B2 => n21165, C1 => n23490, C2 =>
                           n21613, A => n18237, ZN => n18236);
   U15810 : OAI22_X1 port map( A1 => n19553, A2 => n23416, B1 => n19681, B2 => 
                           n23405, ZN => n18238);
   U15811 : AOI221_X1 port map( B1 => n23451, B2 => n21114, C1 => n23435, C2 =>
                           n21543, A => n18184, ZN => n18181);
   U15812 : AOI221_X1 port map( B1 => n23506, B2 => n21185, C1 => n23490, C2 =>
                           n21599, A => n18183, ZN => n18182);
   U15813 : OAI22_X1 port map( A1 => n19554, A2 => n23416, B1 => n19682, B2 => 
                           n23410, ZN => n18184);
   U15814 : AOI221_X1 port map( B1 => n23452, B2 => n21111, C1 => n23436, C2 =>
                           n21540, A => n18400, ZN => n18397);
   U15815 : AOI221_X1 port map( B1 => n23507, B2 => n21183, C1 => n23491, C2 =>
                           n21596, A => n18399, ZN => n18398);
   U15816 : OAI22_X1 port map( A1 => n19550, A2 => n23417, B1 => n19678, B2 => 
                           n23406, ZN => n18400);
   U15817 : AOI221_X1 port map( B1 => n23451, B2 => n21112, C1 => n23435, C2 =>
                           n21541, A => n18346, ZN => n18343);
   U15818 : AOI221_X1 port map( B1 => n23506, B2 => n21184, C1 => n23490, C2 =>
                           n21597, A => n18345, ZN => n18344);
   U15819 : OAI22_X1 port map( A1 => n19551, A2 => n23418, B1 => n19679, B2 => 
                           n23405, ZN => n18346);
   U15820 : AOI221_X1 port map( B1 => n23452, B2 => n21095, C1 => n23436, C2 =>
                           n21524, A => n18373, ZN => n18370);
   U15821 : AOI221_X1 port map( B1 => n23507, B2 => n21174, C1 => n23491, C2 =>
                           n21580, A => n18372, ZN => n18371);
   U15822 : OAI22_X1 port map( A1 => n19545, A2 => n23419, B1 => n19673, B2 => 
                           n23405, ZN => n18373);
   U15823 : AOI221_X1 port map( B1 => n23451, B2 => n21113, C1 => n23435, C2 =>
                           n21542, A => n18211, ZN => n18208);
   U15824 : AOI221_X1 port map( B1 => n23506, B2 => n21159, C1 => n23490, C2 =>
                           n21598, A => n18210, ZN => n18209);
   U15825 : OAI22_X1 port map( A1 => n19542, A2 => n23416, B1 => n19670, B2 => 
                           n23405, ZN => n18211);
   U15826 : AOI221_X1 port map( B1 => n23451, B2 => n21126, C1 => n23435, C2 =>
                           n21555, A => n18319, ZN => n18316);
   U15827 : AOI221_X1 port map( B1 => n23506, B2 => n21164, C1 => n23490, C2 =>
                           n21611, A => n18318, ZN => n18317);
   U15828 : OAI22_X1 port map( A1 => n19544, A2 => n23418, B1 => n19672, B2 => 
                           n23405, ZN => n18319);
   U15829 : AOI221_X1 port map( B1 => n23452, B2 => n21109, C1 => n23436, C2 =>
                           n21538, A => n18454, ZN => n18451);
   U15830 : AOI221_X1 port map( B1 => n23507, B2 => n21182, C1 => n23491, C2 =>
                           n21594, A => n18453, ZN => n18452);
   U15831 : OAI22_X1 port map( A1 => n19549, A2 => n23421, B1 => n19677, B2 => 
                           n23408, ZN => n18454);
   U15832 : AOI221_X1 port map( B1 => n23451, B2 => n21150, C1 => n23435, C2 =>
                           n21631, A => n18265, ZN => n18262);
   U15833 : AOI221_X1 port map( B1 => n23506, B2 => n21207, C1 => n23490, C2 =>
                           n21636, A => n18264, ZN => n18263);
   U15834 : OAI22_X1 port map( A1 => n19543, A2 => n23421, B1 => n19671, B2 => 
                           n23405, ZN => n18265);
   U15835 : AOI221_X1 port map( B1 => n23451, B2 => n21127, C1 => n23435, C2 =>
                           n21556, A => n18292, ZN => n18289);
   U15836 : AOI221_X1 port map( B1 => n23506, B2 => n21193, C1 => n23490, C2 =>
                           n21612, A => n18291, ZN => n18290);
   U15837 : OAI22_X1 port map( A1 => n19552, A2 => n23419, B1 => n19680, B2 => 
                           n23405, ZN => n18292);
   U15838 : OAI22_X1 port map( A1 => n19477, A2 => n23475, B1 => n19605, B2 => 
                           n23459, ZN => n18156);
   U15839 : OAI22_X1 port map( A1 => n19475, A2 => n23473, B1 => n19603, B2 => 
                           n23460, ZN => n18048);
   U15840 : OAI22_X1 port map( A1 => n19492, A2 => n23471, B1 => n19620, B2 => 
                           n23464, ZN => n18075);
   U15841 : AOI221_X1 port map( B1 => n23450, B2 => n21129, C1 => n23434, C2 =>
                           n21558, A => n18157, ZN => n18154);
   U15842 : AOI221_X1 port map( B1 => n23505, B2 => n21194, C1 => n23489, C2 =>
                           n21614, A => n18156, ZN => n18155);
   U15843 : OAI22_X1 port map( A1 => n19541, A2 => n23416, B1 => n19669, B2 => 
                           n23405, ZN => n18157);
   U15844 : AOI221_X1 port map( B1 => n23450, B2 => n21130, C1 => n23434, C2 =>
                           n21559, A => n18049, ZN => n18046);
   U15845 : AOI221_X1 port map( B1 => n23505, B2 => n21166, C1 => n23489, C2 =>
                           n21615, A => n18048, ZN => n18047);
   U15846 : OAI22_X1 port map( A1 => n19539, A2 => n23416, B1 => n19667, B2 => 
                           n23405, ZN => n18049);
   U15847 : AOI221_X1 port map( B1 => n23450, B2 => n21116, C1 => n23434, C2 =>
                           n21545, A => n18076, ZN => n18073);
   U15848 : AOI221_X1 port map( B1 => n23505, B2 => n21187, C1 => n23489, C2 =>
                           n21601, A => n18075, ZN => n18074);
   U15849 : OAI22_X1 port map( A1 => n19556, A2 => n23416, B1 => n19684, B2 => 
                           n23410, ZN => n18076);
   U15850 : OAI22_X1 port map( A1 => n19491, A2 => n23471, B1 => n19619, B2 => 
                           n23464, ZN => n18129);
   U15851 : OAI22_X1 port map( A1 => n19476, A2 => n23474, B1 => n19604, B2 => 
                           n23462, ZN => n18102);
   U15852 : AOI221_X1 port map( B1 => n23450, B2 => n21115, C1 => n23434, C2 =>
                           n21544, A => n18130, ZN => n18127);
   U15853 : AOI221_X1 port map( B1 => n23505, B2 => n21186, C1 => n23489, C2 =>
                           n21600, A => n18129, ZN => n18128);
   U15854 : OAI22_X1 port map( A1 => n19555, A2 => n23416, B1 => n19683, B2 => 
                           n23410, ZN => n18130);
   U15855 : AOI221_X1 port map( B1 => n23450, B2 => n21267, C1 => n23434, C2 =>
                           n21752, A => n18103, ZN => n18100);
   U15856 : AOI221_X1 port map( B1 => n23505, B2 => n21278, C1 => n23489, C2 =>
                           n21758, A => n18102, ZN => n18101);
   U15857 : OAI22_X1 port map( A1 => n19540, A2 => n23416, B1 => n19668, B2 => 
                           n23408, ZN => n18103);
   U15858 : BUF_X1 port map( A => n15182, Z => n23907);
   U15859 : NOR3_X1 port map( A1 => n16529, A2 => ADD_RD2(2), A3 => n16580, ZN 
                           => n15182);
   U15860 : OAI22_X1 port map( A1 => n18971, A2 => n23471, B1 => n19099, B2 => 
                           n23459, ZN => n18476);
   U15861 : OAI22_X1 port map( A1 => n18970, A2 => n23471, B1 => n19098, B2 => 
                           n23459, ZN => n18422);
   U15862 : OAI22_X1 port map( A1 => n18977, A2 => n23471, B1 => n19105, B2 => 
                           n23460, ZN => n18233);
   U15863 : OAI22_X1 port map( A1 => n18978, A2 => n23474, B1 => n19106, B2 => 
                           n23459, ZN => n18179);
   U15864 : OAI22_X1 port map( A1 => n18974, A2 => n23471, B1 => n19102, B2 => 
                           n23459, ZN => n18395);
   U15865 : OAI22_X1 port map( A1 => n18975, A2 => n23475, B1 => n19103, B2 => 
                           n23460, ZN => n18341);
   U15866 : OAI22_X1 port map( A1 => n18969, A2 => n23471, B1 => n19097, B2 => 
                           n23459, ZN => n18368);
   U15867 : OAI22_X1 port map( A1 => n18966, A2 => n23474, B1 => n19094, B2 => 
                           n23460, ZN => n18206);
   U15868 : OAI22_X1 port map( A1 => n18968, A2 => n23472, B1 => n19096, B2 => 
                           n23460, ZN => n18314);
   U15869 : OAI22_X1 port map( A1 => n18973, A2 => n23471, B1 => n19101, B2 => 
                           n23459, ZN => n18449);
   U15870 : OAI22_X1 port map( A1 => n18967, A2 => n23475, B1 => n19095, B2 => 
                           n23460, ZN => n18260);
   U15871 : OAI22_X1 port map( A1 => n18976, A2 => n23475, B1 => n19104, B2 => 
                           n23460, ZN => n18287);
   U15872 : AOI221_X1 port map( B1 => n23452, B2 => n20900, C1 => n23436, C2 =>
                           n21640, A => n18477, ZN => n18474);
   U15873 : AOI221_X1 port map( B1 => n23507, B2 => n21210, C1 => n23491, C2 =>
                           n21695, A => n18476, ZN => n18475);
   U15874 : OAI22_X1 port map( A1 => n19035, A2 => n23417, B1 => n19163, B2 => 
                           n23406, ZN => n18477);
   U15875 : AOI221_X1 port map( B1 => n23452, B2 => n20915, C1 => n23436, C2 =>
                           n21655, A => n18423, ZN => n18420);
   U15876 : AOI221_X1 port map( B1 => n23507, B2 => n21226, C1 => n23491, C2 =>
                           n21711, A => n18422, ZN => n18421);
   U15877 : OAI22_X1 port map( A1 => n19034, A2 => n23418, B1 => n19162, B2 => 
                           n23408, ZN => n18423);
   U15878 : AOI221_X1 port map( B1 => n23451, B2 => n20934, C1 => n23435, C2 =>
                           n21674, A => n18234, ZN => n18231);
   U15879 : AOI221_X1 port map( B1 => n23506, B2 => n21246, C1 => n23490, C2 =>
                           n21730, A => n18233, ZN => n18232);
   U15880 : OAI22_X1 port map( A1 => n19041, A2 => n23417, B1 => n19169, B2 => 
                           n23405, ZN => n18234);
   U15881 : AOI221_X1 port map( B1 => n23450, B2 => n20919, C1 => n23434, C2 =>
                           n21659, A => n18180, ZN => n18177);
   U15882 : AOI221_X1 port map( B1 => n23505, B2 => n21230, C1 => n23489, C2 =>
                           n21715, A => n18179, ZN => n18178);
   U15883 : OAI22_X1 port map( A1 => n19042, A2 => n23416, B1 => n19170, B2 => 
                           n23410, ZN => n18180);
   U15884 : AOI221_X1 port map( B1 => n23452, B2 => n20916, C1 => n23436, C2 =>
                           n21656, A => n18396, ZN => n18393);
   U15885 : AOI221_X1 port map( B1 => n23507, B2 => n21227, C1 => n23491, C2 =>
                           n21712, A => n18395, ZN => n18394);
   U15886 : OAI22_X1 port map( A1 => n19038, A2 => n23421, B1 => n19166, B2 => 
                           n23409, ZN => n18396);
   U15887 : AOI221_X1 port map( B1 => n23451, B2 => n20917, C1 => n23435, C2 =>
                           n21657, A => n18342, ZN => n18339);
   U15888 : AOI221_X1 port map( B1 => n23506, B2 => n21228, C1 => n23490, C2 =>
                           n21713, A => n18341, ZN => n18340);
   U15889 : OAI22_X1 port map( A1 => n19039, A2 => n23416, B1 => n19167, B2 => 
                           n23405, ZN => n18342);
   U15890 : AOI221_X1 port map( B1 => n23452, B2 => n20901, C1 => n23436, C2 =>
                           n21641, A => n18369, ZN => n18366);
   U15891 : AOI221_X1 port map( B1 => n23507, B2 => n21211, C1 => n23491, C2 =>
                           n21696, A => n18368, ZN => n18367);
   U15892 : OAI22_X1 port map( A1 => n19033, A2 => n23420, B1 => n19161, B2 => 
                           n23409, ZN => n18369);
   U15893 : AOI221_X1 port map( B1 => n23451, B2 => n20918, C1 => n23435, C2 =>
                           n21658, A => n18207, ZN => n18204);
   U15894 : AOI221_X1 port map( B1 => n23506, B2 => n21229, C1 => n23490, C2 =>
                           n21714, A => n18206, ZN => n18205);
   U15895 : OAI22_X1 port map( A1 => n19030, A2 => n23416, B1 => n19158, B2 => 
                           n23405, ZN => n18207);
   U15896 : AOI221_X1 port map( B1 => n23451, B2 => n20932, C1 => n23435, C2 =>
                           n21672, A => n18315, ZN => n18312);
   U15897 : AOI221_X1 port map( B1 => n23506, B2 => n21244, C1 => n23490, C2 =>
                           n21728, A => n18314, ZN => n18313);
   U15898 : OAI22_X1 port map( A1 => n19032, A2 => n23418, B1 => n19160, B2 => 
                           n23405, ZN => n18315);
   U15899 : AOI221_X1 port map( B1 => n23452, B2 => n20914, C1 => n23436, C2 =>
                           n21654, A => n18450, ZN => n18447);
   U15900 : AOI221_X1 port map( B1 => n23507, B2 => n21225, C1 => n23491, C2 =>
                           n21710, A => n18449, ZN => n18448);
   U15901 : OAI22_X1 port map( A1 => n19037, A2 => n23417, B1 => n19165, B2 => 
                           n23410, ZN => n18450);
   U15902 : AOI221_X1 port map( B1 => n23451, B2 => n20955, C1 => n23435, C2 =>
                           n21751, A => n18261, ZN => n18258);
   U15903 : AOI221_X1 port map( B1 => n23506, B2 => n21266, C1 => n23490, C2 =>
                           n21754, A => n18260, ZN => n18259);
   U15904 : OAI22_X1 port map( A1 => n19031, A2 => n23420, B1 => n19159, B2 => 
                           n23405, ZN => n18261);
   U15905 : AOI221_X1 port map( B1 => n23451, B2 => n20933, C1 => n23435, C2 =>
                           n21673, A => n18288, ZN => n18285);
   U15906 : AOI221_X1 port map( B1 => n23506, B2 => n21245, C1 => n23490, C2 =>
                           n21729, A => n18287, ZN => n18286);
   U15907 : OAI22_X1 port map( A1 => n19040, A2 => n23419, B1 => n19168, B2 => 
                           n23405, ZN => n18288);
   U15908 : OAI22_X1 port map( A1 => n18979, A2 => n23471, B1 => n19107, B2 => 
                           n23460, ZN => n18125);
   U15909 : OAI22_X1 port map( A1 => n18965, A2 => n23474, B1 => n19093, B2 => 
                           n23461, ZN => n18152);
   U15910 : OAI22_X1 port map( A1 => n18964, A2 => n23471, B1 => n19092, B2 => 
                           n23464, ZN => n18098);
   U15911 : OAI22_X1 port map( A1 => n18963, A2 => n23473, B1 => n19091, B2 => 
                           n23463, ZN => n18044);
   U15912 : OAI22_X1 port map( A1 => n18980, A2 => n23473, B1 => n19108, B2 => 
                           n23464, ZN => n18071);
   U15913 : AOI221_X1 port map( B1 => n23450, B2 => n20920, C1 => n23434, C2 =>
                           n21660, A => n18126, ZN => n18123);
   U15914 : AOI221_X1 port map( B1 => n23505, B2 => n21231, C1 => n23489, C2 =>
                           n21716, A => n18125, ZN => n18124);
   U15915 : OAI22_X1 port map( A1 => n19043, A2 => n23416, B1 => n19171, B2 => 
                           n23405, ZN => n18126);
   U15916 : AOI221_X1 port map( B1 => n23450, B2 => n20935, C1 => n23434, C2 =>
                           n21675, A => n18153, ZN => n18150);
   U15917 : AOI221_X1 port map( B1 => n23505, B2 => n21247, C1 => n23489, C2 =>
                           n21731, A => n18152, ZN => n18151);
   U15918 : OAI22_X1 port map( A1 => n19029, A2 => n23416, B1 => n19157, B2 => 
                           n23406, ZN => n18153);
   U15919 : AOI221_X1 port map( B1 => n23450, B2 => n20957, C1 => n23434, C2 =>
                           n21830, A => n18099, ZN => n18096);
   U15920 : AOI221_X1 port map( B1 => n23505, B2 => n21279, C1 => n23489, C2 =>
                           n21835, A => n18098, ZN => n18097);
   U15921 : OAI22_X1 port map( A1 => n19028, A2 => n23416, B1 => n19156, B2 => 
                           n23407, ZN => n18099);
   U15922 : AOI221_X1 port map( B1 => n23450, B2 => n20936, C1 => n23434, C2 =>
                           n21676, A => n18045, ZN => n18042);
   U15923 : AOI221_X1 port map( B1 => n23505, B2 => n21248, C1 => n23489, C2 =>
                           n21732, A => n18044, ZN => n18043);
   U15924 : OAI22_X1 port map( A1 => n19027, A2 => n23416, B1 => n19155, B2 => 
                           n23408, ZN => n18045);
   U15925 : AOI221_X1 port map( B1 => n23450, B2 => n20921, C1 => n23434, C2 =>
                           n21661, A => n18072, ZN => n18069);
   U15926 : AOI221_X1 port map( B1 => n23505, B2 => n21232, C1 => n23489, C2 =>
                           n21717, A => n18071, ZN => n18070);
   U15927 : OAI22_X1 port map( A1 => n19044, A2 => n23416, B1 => n19172, B2 => 
                           n23410, ZN => n18072);
   U15928 : OAI22_X1 port map( A1 => n19484, A2 => n23471, B1 => n19612, B2 => 
                           n23459, ZN => n18519);
   U15929 : AOI221_X1 port map( B1 => n23452, B2 => n21284, C1 => n23436, C2 =>
                           n21841, A => n18520, ZN => n18517);
   U15930 : AOI221_X1 port map( B1 => n23507, B2 => n21286, C1 => n23491, C2 =>
                           n21840, A => n18519, ZN => n18518);
   U15931 : OAI22_X1 port map( A1 => n19548, A2 => n23421, B1 => n19676, B2 => 
                           n23407, ZN => n18520);
   U15932 : OAI22_X1 port map( A1 => n18972, A2 => n23471, B1 => n19100, B2 => 
                           n23459, ZN => n18515);
   U15933 : AOI221_X1 port map( B1 => n23452, B2 => n20962, C1 => n23436, C2 =>
                           n21843, A => n18516, ZN => n18513);
   U15934 : AOI221_X1 port map( B1 => n23507, B2 => n21285, C1 => n23491, C2 =>
                           n21842, A => n18515, ZN => n18514);
   U15935 : OAI22_X1 port map( A1 => n19036, A2 => n23416, B1 => n19164, B2 => 
                           n23406, ZN => n18516);
   U15936 : BUF_X1 port map( A => n15183, Z => n23898);
   U15937 : NOR3_X1 port map( A1 => n16579, A2 => RESET, A3 => n23946, ZN => 
                           n15183);
   U15938 : NOR3_X1 port map( A1 => n25404, A2 => ADD_WR(0), A3 => n16668, ZN 
                           => n16678);
   U15939 : NOR3_X1 port map( A1 => n16668, A2 => ADD_WR(1), A3 => n25405, ZN 
                           => n16673);
   U15940 : AOI21_X1 port map( B1 => n16580, B2 => ADD_RD2(2), A => ADD_RD2(3),
                           ZN => n16579);
   U15941 : INV_X1 port map( A => ADD_RD1(2), ZN => n24369);
   U15942 : AND2_X1 port map( A1 => SIGRETURN, A2 => n23037, ZN => n22767);
   U15943 : INV_X1 port map( A => ADD_RD2(1), ZN => n25408);
   U15944 : INV_X1 port map( A => ADD_RD2(0), ZN => n25409);
   U15945 : CLKBUF_X1 port map( A => n23014, Z => n22769);
   U15946 : BUF_X2 port map( A => n22489, Z => n23014);
   U15947 : BUF_X1 port map( A => n23015, Z => n22771);
   U15948 : INV_X1 port map( A => n24090, ZN => n22772);
   U15949 : INV_X1 port map( A => n22772, ZN => n22773);
   U15950 : INV_X1 port map( A => n22772, ZN => n22774);
   U15951 : INV_X1 port map( A => n22772, ZN => n22775);
   U15952 : INV_X1 port map( A => n22776, ZN => n22777);
   U15953 : INV_X1 port map( A => n22776, ZN => n22778);
   U15954 : INV_X1 port map( A => n22776, ZN => n22779);
   U15955 : CLKBUF_X1 port map( A => n24183, Z => n22796);
   U15956 : CLKBUF_X1 port map( A => n24183, Z => n22797);
   U15957 : CLKBUF_X2 port map( A => n25379, Z => n22798);
   U15958 : BUF_X4 port map( A => n25379, Z => n22799);
   U15959 : CLKBUF_X2 port map( A => n25379, Z => n22800);
   U15960 : NAND2_X1 port map( A1 => n21456, A2 => n24358, ZN => n25379);
   U15961 : INV_X1 port map( A => n24349, ZN => n22802);
   U15962 : BUF_X1 port map( A => n22802, Z => n22803);
   U15963 : BUF_X1 port map( A => n22802, Z => n22804);
   U15964 : BUF_X1 port map( A => n22802, Z => n22805);
   U15965 : BUF_X1 port map( A => n22802, Z => n22806);
   U15966 : BUF_X1 port map( A => n22802, Z => n22807);
   U15967 : BUF_X1 port map( A => n22802, Z => n22808);
   U15968 : BUF_X1 port map( A => n22802, Z => n22809);
   U15969 : BUF_X1 port map( A => n22802, Z => n22810);
   U15970 : BUF_X1 port map( A => n22802, Z => n22811);
   U15971 : BUF_X1 port map( A => n22802, Z => n22812);
   U15972 : INV_X1 port map( A => n22798, ZN => n22909);
   U15973 : INV_X1 port map( A => n24345, ZN => n22910);
   U15974 : BUF_X1 port map( A => n22910, Z => n22919);
   U15975 : BUF_X1 port map( A => n22910, Z => n22920);
   U15976 : BUF_X2 port map( A => n25383, Z => n22922);
   U15977 : BUF_X2 port map( A => n25383, Z => n22923);
   U15978 : INV_X1 port map( A => n24376, ZN => n25383);
   U15979 : AND2_X1 port map( A1 => n22918, A2 => n22199, ZN => n22924);
   U15980 : AND2_X1 port map( A1 => n22805, A2 => n21278, ZN => n22925);
   U15981 : NOR3_X1 port map( A1 => n22924, A2 => n22925, A3 => n24611, ZN => 
                           n24617);
   U15982 : AND2_X1 port map( A1 => n22919, A2 => n22198, ZN => n22926);
   U15983 : AND2_X1 port map( A1 => n22802, A2 => n21186, ZN => n22927);
   U15984 : NOR3_X1 port map( A1 => n22926, A2 => n22927, A3 => n24595, ZN => 
                           n24601);
   U15985 : AND2_X1 port map( A1 => n22923, A2 => n22188, ZN => n22928);
   U15986 : AND2_X1 port map( A1 => n22969, A2 => n21271, ZN => n22929);
   U15987 : NOR3_X1 port map( A1 => n22928, A2 => n22929, A3 => n24962, ZN => 
                           n24970);
   U15988 : AND2_X1 port map( A1 => n22523, A2 => n22224, ZN => n22938);
   U15989 : AND2_X1 port map( A1 => n22971, A2 => n21208, ZN => n22939);
   U15990 : NOR3_X1 port map( A1 => n22938, A2 => n22939, A3 => n24722, ZN => 
                           n24730);
   U15991 : OR2_X1 port map( A1 => n19559, A2 => n22934, ZN => n22940);
   U15992 : OR2_X1 port map( A1 => n24721, A2 => n22798, ZN => n22941);
   U15993 : OR2_X1 port map( A1 => n19687, A2 => n22521, ZN => n22942);
   U15994 : NAND3_X1 port map( A1 => n22940, A2 => n22941, A3 => n22942, ZN => 
                           n24722);
   U15995 : BUF_X2 port map( A => n22969, Z => n22971);
   U15996 : AOI221_X1 port map( B1 => n23277, B2 => n20899, C1 => n22494, C2 =>
                           n21639, A => n24758, ZN => n24759);
   U15997 : INV_X1 port map( A => n22633, ZN => n23268);
   U15998 : INV_X1 port map( A => n24354, ZN => n22956);
   U15999 : BUF_X1 port map( A => n22956, Z => n22958);
   U16000 : BUF_X1 port map( A => n22956, Z => n22959);
   U16001 : BUF_X1 port map( A => n22956, Z => n22960);
   U16002 : BUF_X1 port map( A => n22956, Z => n22961);
   U16003 : INV_X1 port map( A => n24354, ZN => n22962);
   U16004 : INV_X1 port map( A => n24386, ZN => n22963);
   U16005 : BUF_X1 port map( A => n25388, Z => n22968);
   U16006 : INV_X4 port map( A => n24386, ZN => n25391);
   U16007 : INV_X1 port map( A => n24344, ZN => n22969);
   U16008 : BUF_X1 port map( A => n22969, Z => n22970);
   U16009 : BUF_X1 port map( A => n22969, Z => n22972);
   U16010 : BUF_X1 port map( A => n22969, Z => n22973);
   U16011 : BUF_X1 port map( A => n22969, Z => n22974);
   U16012 : INV_X1 port map( A => n24344, ZN => n22975);
   U16013 : BUF_X2 port map( A => n23010, Z => n23009);
   U16014 : INV_X1 port map( A => RESET, ZN => n25403);
   U16015 : INV_X1 port map( A => CALL, ZN => n24127);
   U16016 : INV_X1 port map( A => SIGRETURN, ZN => n24002);
   U16017 : NAND2_X1 port map( A1 => n23037, A2 => n24002, ZN => n24010);
   U16018 : INV_X1 port map( A => n24010, ZN => n24342);
   U16019 : OAI21_X1 port map( B1 => n22690, B2 => n23053, A => n24342, ZN => 
                           n23981);
   U16020 : INV_X1 port map( A => n3259, ZN => n24143);
   U16021 : NAND2_X1 port map( A1 => n23948, A2 => n22499, ZN => n24341);
   U16022 : NAND2_X1 port map( A1 => n22988, A2 => n22493, ZN => n23949);
   U16023 : OAI22_X1 port map( A1 => i_0_port, A2 => n23949, B1 => n3242, B2 =>
                           n22988, ZN => n13242);
   U16024 : INV_X1 port map( A => n23949, ZN => n23980);
   U16025 : AOI22_X1 port map( A1 => n22987, A2 => i_31_port, B1 => N653, B2 =>
                           n22984, ZN => n23950);
   U16026 : INV_X1 port map( A => n23950, ZN => n13211);
   U16027 : AOI22_X1 port map( A1 => n22987, A2 => i_30_port, B1 => N652, B2 =>
                           n22984, ZN => n23951);
   U16028 : INV_X1 port map( A => n23951, ZN => n13212);
   U16029 : AOI22_X1 port map( A1 => n22987, A2 => i_29_port, B1 => N651, B2 =>
                           n22984, ZN => n23952);
   U16030 : INV_X1 port map( A => n23952, ZN => n13213);
   U16031 : AOI22_X1 port map( A1 => n22987, A2 => i_28_port, B1 => N650, B2 =>
                           n22984, ZN => n23953);
   U16032 : INV_X1 port map( A => n23953, ZN => n13214);
   U16033 : AOI22_X1 port map( A1 => n22987, A2 => i_27_port, B1 => N649, B2 =>
                           n22984, ZN => n23954);
   U16034 : INV_X1 port map( A => n23954, ZN => n13215);
   U16035 : AOI22_X1 port map( A1 => n22987, A2 => i_26_port, B1 => N648, B2 =>
                           n22984, ZN => n23955);
   U16036 : INV_X1 port map( A => n23955, ZN => n13216);
   U16037 : AOI22_X1 port map( A1 => n22987, A2 => i_25_port, B1 => N647, B2 =>
                           n22984, ZN => n23956);
   U16038 : INV_X1 port map( A => n23956, ZN => n13217);
   U16039 : AOI22_X1 port map( A1 => n22987, A2 => i_24_port, B1 => N646, B2 =>
                           n22984, ZN => n23957);
   U16040 : INV_X1 port map( A => n23957, ZN => n13218);
   U16041 : AOI22_X1 port map( A1 => n22987, A2 => i_23_port, B1 => N645, B2 =>
                           n22984, ZN => n23958);
   U16042 : INV_X1 port map( A => n23958, ZN => n13219);
   U16043 : AOI22_X1 port map( A1 => n22987, A2 => i_22_port, B1 => N644, B2 =>
                           n22984, ZN => n23959);
   U16044 : INV_X1 port map( A => n23959, ZN => n13220);
   U16045 : AOI22_X1 port map( A1 => n22987, A2 => i_21_port, B1 => N643, B2 =>
                           n22984, ZN => n23960);
   U16046 : INV_X1 port map( A => n23960, ZN => n13221);
   U16047 : AOI22_X1 port map( A1 => n22987, A2 => i_20_port, B1 => N642, B2 =>
                           n22984, ZN => n23961);
   U16048 : INV_X1 port map( A => n23961, ZN => n13222);
   U16049 : AOI22_X1 port map( A1 => n23981, A2 => i_19_port, B1 => N641, B2 =>
                           n22985, ZN => n23962);
   U16050 : INV_X1 port map( A => n23962, ZN => n13223);
   U16051 : AOI22_X1 port map( A1 => n23981, A2 => i_18_port, B1 => N640, B2 =>
                           n22985, ZN => n23963);
   U16052 : INV_X1 port map( A => n23963, ZN => n13224);
   U16053 : AOI22_X1 port map( A1 => n23981, A2 => i_17_port, B1 => N639, B2 =>
                           n22985, ZN => n23964);
   U16054 : INV_X1 port map( A => n23964, ZN => n13225);
   U16055 : AOI22_X1 port map( A1 => n22987, A2 => i_16_port, B1 => N638, B2 =>
                           n22985, ZN => n23965);
   U16056 : INV_X1 port map( A => n23965, ZN => n13226);
   U16057 : AOI22_X1 port map( A1 => n22987, A2 => i_15_port, B1 => N637, B2 =>
                           n22985, ZN => n23966);
   U16058 : INV_X1 port map( A => n23966, ZN => n13227);
   U16059 : AOI22_X1 port map( A1 => n22987, A2 => i_14_port, B1 => N636, B2 =>
                           n22985, ZN => n23967);
   U16060 : INV_X1 port map( A => n23967, ZN => n13228);
   U16061 : AOI22_X1 port map( A1 => n22987, A2 => i_13_port, B1 => N635, B2 =>
                           n22985, ZN => n23968);
   U16062 : INV_X1 port map( A => n23968, ZN => n13229);
   U16063 : AOI22_X1 port map( A1 => n22987, A2 => i_12_port, B1 => N634, B2 =>
                           n22985, ZN => n23969);
   U16064 : INV_X1 port map( A => n23969, ZN => n13230);
   U16065 : AOI22_X1 port map( A1 => n22987, A2 => i_11_port, B1 => N633, B2 =>
                           n22985, ZN => n23970);
   U16066 : INV_X1 port map( A => n23970, ZN => n13231);
   U16067 : AOI22_X1 port map( A1 => n22987, A2 => i_10_port, B1 => N632, B2 =>
                           n22985, ZN => n23971);
   U16068 : INV_X1 port map( A => n23971, ZN => n13232);
   U16069 : AOI22_X1 port map( A1 => n22987, A2 => i_9_port, B1 => N631, B2 => 
                           n22985, ZN => n23972);
   U16070 : INV_X1 port map( A => n23972, ZN => n13233);
   U16071 : AOI22_X1 port map( A1 => n22987, A2 => i_8_port, B1 => N630, B2 => 
                           n22985, ZN => n23973);
   U16072 : INV_X1 port map( A => n23973, ZN => n13234);
   U16073 : AOI22_X1 port map( A1 => n22987, A2 => i_7_port, B1 => N629, B2 => 
                           n22986, ZN => n23974);
   U16074 : INV_X1 port map( A => n23974, ZN => n13235);
   U16075 : AOI22_X1 port map( A1 => n23981, A2 => i_6_port, B1 => N628, B2 => 
                           n22986, ZN => n23975);
   U16076 : INV_X1 port map( A => n23975, ZN => n13236);
   U16077 : AOI22_X1 port map( A1 => n22987, A2 => i_5_port, B1 => N627, B2 => 
                           n22986, ZN => n23976);
   U16078 : INV_X1 port map( A => n23976, ZN => n13237);
   U16079 : AOI22_X1 port map( A1 => n23981, A2 => i_4_port, B1 => N626, B2 => 
                           n22986, ZN => n23977);
   U16080 : INV_X1 port map( A => n23977, ZN => n13238);
   U16081 : AOI22_X1 port map( A1 => n22987, A2 => n24143, B1 => N624, B2 => 
                           n22986, ZN => n23978);
   U16082 : INV_X1 port map( A => n23978, ZN => n13240);
   U16083 : AOI22_X1 port map( A1 => n23981, A2 => i_1_port, B1 => N623, B2 => 
                           n22986, ZN => n23979);
   U16084 : INV_X1 port map( A => n23979, ZN => n13241);
   U16085 : AOI22_X1 port map( A1 => n22987, A2 => i_3_port, B1 => N625, B2 => 
                           n22986, ZN => n23982);
   U16086 : INV_X1 port map( A => n23982, ZN => n13239);
   U16087 : NAND3_X1 port map( A1 => n22769, A2 => n23284, A3 => n23037, ZN => 
                           n23984);
   U16088 : INV_X1 port map( A => n23984, ZN => n24338);
   U16089 : NAND2_X1 port map( A1 => CALL, A2 => n23283, ZN => n24337);
   U16090 : OAI21_X1 port map( B1 => n22768, B2 => n23186, A => n24337, ZN => 
                           n5642);
   U16091 : NAND2_X1 port map( A1 => n5699, A2 => n24002, ZN => n24086);
   U16092 : NAND4_X1 port map( A1 => n23053, A2 => n24008, A3 => n22512, A4 => 
                           n23037, ZN => n23983);
   U16093 : INV_X1 port map( A => n23983, ZN => n24340);
   U16094 : NAND2_X1 port map( A1 => n23006, A2 => n23283, ZN => n24339);
   U16095 : OAI21_X1 port map( B1 => n5700, B2 => n24340, A => n24339, ZN => 
                           n5641);
   U16096 : MUX2_X1 port map( A => n21416, B => n22506, S => n23186, Z => n5646
                           );
   U16097 : INV_X1 port map( A => N210, ZN => n24185);
   U16098 : NAND2_X1 port map( A1 => n22768, A2 => n22990, ZN => n24000);
   U16099 : INV_X1 port map( A => n24000, ZN => n23992);
   U16100 : NAND4_X1 port map( A1 => n24073, A2 => n22539, A3 => n22540, A4 => 
                           n22541, ZN => n23988);
   U16101 : NAND4_X1 port map( A1 => n24047, A2 => n24045, A3 => n22780, A4 => 
                           n24065, ZN => n23987);
   U16102 : NAND4_X1 port map( A1 => n22783, A2 => n22785, A3 => n22789, A4 => 
                           n22790, ZN => n23986);
   U16103 : NAND4_X1 port map( A1 => n22786, A2 => n22793, A3 => n22795, A4 => 
                           n22981, ZN => n23985);
   U16104 : NOR4_X1 port map( A1 => n23987, A2 => n23988, A3 => n23986, A4 => 
                           n23985, ZN => n23989);
   U16105 : NAND2_X1 port map( A1 => n23990, A2 => n23989, ZN => n24087);
   U16106 : OAI222_X1 port map( A1 => n5756, A2 => n22997, B1 => n22505, B2 => 
                           n22994, C1 => n22788, C2 => n22990, ZN => n5645);
   U16107 : MUX2_X1 port map( A => n21417, B => n22498, S => n23186, Z => n5609
                           );
   U16108 : INV_X1 port map( A => N211, ZN => n24184);
   U16109 : OAI222_X1 port map( A1 => n5755, A2 => n22997, B1 => n22497, B2 => 
                           n22994, C1 => n22982, C2 => n22991, ZN => n5448);
   U16110 : MUX2_X1 port map( A => n21419, B => n22532, S => n23186, Z => n5610
                           );
   U16111 : INV_X1 port map( A => N212, ZN => n24183);
   U16112 : OAI222_X1 port map( A1 => n5747, A2 => n22997, B1 => n22796, B2 => 
                           n22994, C1 => n22983, C2 => n22991, ZN => n5447);
   U16113 : MUX2_X1 port map( A => n21418, B => n22547, S => n23186, Z => n5611
                           );
   U16114 : INV_X1 port map( A => N213, ZN => n24290);
   U16115 : OAI222_X1 port map( A1 => n5736, A2 => n22997, B1 => n24290, B2 => 
                           n22994, C1 => n22784, C2 => n22991, ZN => n5446);
   U16116 : MUX2_X1 port map( A => n21420, B => n22495, S => n23186, Z => n5612
                           );
   U16117 : INV_X1 port map( A => N214, ZN => n24138);
   U16118 : OAI222_X1 port map( A1 => n5733, A2 => n22997, B1 => n24138, B2 => 
                           n22994, C1 => n22787, C2 => n22991, ZN => n5445);
   U16119 : MUX2_X1 port map( A => n21421, B => n22511, S => n23186, Z => n5614
                           );
   U16120 : INV_X1 port map( A => n22511, ZN => n24123);
   U16121 : OAI222_X1 port map( A1 => n5732, A2 => n22997, B1 => n24123, B2 => 
                           n22994, C1 => n22791, C2 => n22991, ZN => n5444);
   U16122 : MUX2_X1 port map( A => n21424, B => N218, S => n23186, Z => n5616);
   U16123 : INV_X1 port map( A => N218, ZN => n24121);
   U16124 : OAI222_X1 port map( A1 => n5731, A2 => n22997, B1 => n24121, B2 => 
                           n22994, C1 => n22792, C2 => n22991, ZN => n5443);
   U16125 : MUX2_X1 port map( A => n21028, B => N221, S => n23186, Z => n5619);
   U16126 : INV_X1 port map( A => N221, ZN => n24118);
   U16127 : OAI222_X1 port map( A1 => n5754, A2 => n22997, B1 => n24118, B2 => 
                           n22994, C1 => n24071, C2 => n22991, ZN => n5442);
   U16128 : MUX2_X1 port map( A => n21427, B => N222, S => n23185, Z => n5620);
   U16129 : INV_X1 port map( A => N222, ZN => n24117);
   U16130 : OAI222_X1 port map( A1 => n5753, A2 => n22997, B1 => n24117, B2 => 
                           n22994, C1 => n24069, C2 => n22991, ZN => n5441);
   U16131 : MUX2_X1 port map( A => n21426, B => n22530, S => n23185, Z => n5621
                           );
   U16132 : INV_X1 port map( A => N223, ZN => n24116);
   U16133 : OAI222_X1 port map( A1 => n5752, A2 => n22997, B1 => n24116, B2 => 
                           n22994, C1 => n22781, C2 => n22991, ZN => n5440);
   U16134 : MUX2_X1 port map( A => n21029, B => N224, S => n23185, Z => n5622);
   U16135 : INV_X1 port map( A => N224, ZN => n24115);
   U16136 : OAI222_X1 port map( A1 => n5751, A2 => n22997, B1 => n24115, B2 => 
                           n22994, C1 => n22782, C2 => n22991, ZN => n5439);
   U16137 : MUX2_X1 port map( A => n21431, B => N227, S => n23185, Z => n5625);
   U16138 : INV_X1 port map( A => N227, ZN => n24112);
   U16139 : OAI222_X1 port map( A1 => n5750, A2 => n22997, B1 => n24112, B2 => 
                           n22994, C1 => n24062, C2 => n22991, ZN => n5438);
   U16140 : MUX2_X1 port map( A => n21430, B => N228, S => n23185, Z => n5626);
   U16141 : INV_X1 port map( A => N228, ZN => n24111);
   U16142 : OAI222_X1 port map( A1 => n5749, A2 => n22997, B1 => n24111, B2 => 
                           n22995, C1 => n24060, C2 => n22991, ZN => n5437);
   U16143 : MUX2_X1 port map( A => n21030, B => N229, S => n23185, Z => n5627);
   U16144 : INV_X1 port map( A => N229, ZN => n24110);
   U16145 : OAI222_X1 port map( A1 => n5748, A2 => n22997, B1 => n22500, B2 => 
                           n22995, C1 => n24058, C2 => n22991, ZN => n5436);
   U16146 : MUX2_X1 port map( A => n21435, B => N230, S => n23185, Z => n5628);
   U16147 : INV_X1 port map( A => N230, ZN => n24109);
   U16148 : OAI222_X1 port map( A1 => n5746, A2 => n22997, B1 => n24109, B2 => 
                           n22995, C1 => n22509, C2 => n22991, ZN => n5435);
   U16149 : MUX2_X1 port map( A => n21436, B => N231, S => n23185, Z => n5629);
   U16150 : INV_X1 port map( A => N231, ZN => n24108);
   U16151 : OAI222_X1 port map( A1 => n5745, A2 => n22997, B1 => n24108, B2 => 
                           n22995, C1 => n22786, C2 => n22991, ZN => n5434);
   U16152 : MUX2_X1 port map( A => n21433, B => N232, S => n23185, Z => n5630);
   U16153 : INV_X1 port map( A => N232, ZN => n24107);
   U16154 : OAI222_X1 port map( A1 => n5744, A2 => n22997, B1 => n24107, B2 => 
                           n22995, C1 => n22793, C2 => n22990, ZN => n5433);
   U16155 : MUX2_X1 port map( A => n21434, B => N233, S => n23185, Z => n5631);
   U16156 : INV_X1 port map( A => N233, ZN => n24106);
   U16157 : OAI222_X1 port map( A1 => n5743, A2 => n22997, B1 => n24106, B2 => 
                           n22995, C1 => n22795, C2 => n22990, ZN => n5432);
   U16158 : MUX2_X1 port map( A => n21437, B => N234, S => n23185, Z => n5632);
   U16159 : INV_X1 port map( A => N234, ZN => n24105);
   U16160 : OAI222_X1 port map( A1 => n5742, A2 => n22997, B1 => n24105, B2 => 
                           n22995, C1 => n22981, C2 => n22990, ZN => n5431);
   U16161 : MUX2_X1 port map( A => n21439, B => N235, S => n23184, Z => n5633);
   U16162 : INV_X1 port map( A => N235, ZN => n24104);
   U16163 : OAI222_X1 port map( A1 => n5741, A2 => n22997, B1 => n24104, B2 => 
                           n22995, C1 => n22783, C2 => n22990, ZN => n5430);
   U16164 : MUX2_X1 port map( A => n21441, B => N236, S => n23184, Z => n5634);
   U16165 : INV_X1 port map( A => N236, ZN => n24103);
   U16166 : OAI222_X1 port map( A1 => n5740, A2 => n22997, B1 => n24103, B2 => 
                           n22995, C1 => n22785, C2 => n22990, ZN => n5429);
   U16167 : MUX2_X1 port map( A => n21442, B => N237, S => n23184, Z => n5635);
   U16168 : INV_X1 port map( A => N237, ZN => n24102);
   U16169 : OAI222_X1 port map( A1 => n5739, A2 => n22997, B1 => n24102, B2 => 
                           n22995, C1 => n22789, C2 => n22990, ZN => n5428);
   U16170 : MUX2_X1 port map( A => n21446, B => N238, S => n23184, Z => n5636);
   U16171 : INV_X1 port map( A => N238, ZN => n24101);
   U16172 : OAI222_X1 port map( A1 => n5738, A2 => n22997, B1 => n24101, B2 => 
                           n22995, C1 => n22790, C2 => n22990, ZN => n5427);
   U16173 : MUX2_X1 port map( A => n21449, B => N239, S => n23184, Z => n5637);
   U16174 : INV_X1 port map( A => N239, ZN => n24100);
   U16175 : OAI222_X1 port map( A1 => n5737, A2 => n22997, B1 => n24100, B2 => 
                           n22995, C1 => n24047, C2 => n22990, ZN => n5426);
   U16176 : MUX2_X1 port map( A => n21453, B => N240, S => n23185, Z => n5638);
   U16177 : INV_X1 port map( A => N240, ZN => n24099);
   U16178 : OAI222_X1 port map( A1 => n5735, A2 => n22997, B1 => n24099, B2 => 
                           n22996, C1 => n24045, C2 => n22990, ZN => n5425);
   U16179 : MUX2_X1 port map( A => n21432, B => N226, S => n23184, Z => n5624);
   U16180 : INV_X1 port map( A => n22510, ZN => n23991);
   U16181 : NAND2_X1 port map( A1 => n23991, A2 => n23992, ZN => n23999);
   U16182 : AOI22_X1 port map( A1 => n23992, A2 => N226, B1 => n22999, B2 => 
                           n21432, ZN => n23993);
   U16183 : OAI211_X1 port map( C1 => n22780, C2 => n22991, A => n23999, B => 
                           n23993, ZN => n5424);
   U16184 : MUX2_X1 port map( A => n21428, B => n22513, S => n23184, Z => n5623
                           );
   U16185 : INV_X1 port map( A => n22513, ZN => n24114);
   U16186 : AOI22_X1 port map( A1 => n22999, A2 => n21428, B1 => n22993, B2 => 
                           n20756, ZN => n23994);
   U16187 : OAI211_X1 port map( C1 => n24114, C2 => n24000, A => n23999, B => 
                           n23994, ZN => n5423);
   U16188 : MUX2_X1 port map( A => n21425, B => n22528, S => n23184, Z => n5618
                           );
   U16189 : INV_X1 port map( A => N220, ZN => n24119);
   U16190 : AOI22_X1 port map( A1 => n22999, A2 => n21425, B1 => n22993, B2 => 
                           n20761, ZN => n23995);
   U16191 : OAI211_X1 port map( C1 => n22504, C2 => n24000, A => n23999, B => 
                           n23995, ZN => n5422);
   U16192 : MUX2_X1 port map( A => n21027, B => N219, S => n23184, Z => n5617);
   U16193 : INV_X1 port map( A => N219, ZN => n24120);
   U16194 : AOI22_X1 port map( A1 => n22999, A2 => n21027, B1 => n22993, B2 => 
                           n20732, ZN => n23996);
   U16195 : OAI211_X1 port map( C1 => n22531, C2 => n24000, A => n23999, B => 
                           n23996, ZN => n5421);
   U16196 : MUX2_X1 port map( A => n21423, B => n22503, S => n23184, Z => n5615
                           );
   U16197 : INV_X1 port map( A => n22503, ZN => n24122);
   U16198 : AOI22_X1 port map( A1 => n22999, A2 => n21423, B1 => n22993, B2 => 
                           n20734, ZN => n23997);
   U16199 : OAI211_X1 port map( C1 => n24122, C2 => n24000, A => n23999, B => 
                           n23997, ZN => n5420);
   U16200 : MUX2_X1 port map( A => n21422, B => n22542, S => n23184, Z => n5613
                           );
   U16201 : INV_X1 port map( A => N215, ZN => n24124);
   U16202 : AOI22_X1 port map( A1 => n22999, A2 => n21422, B1 => n22993, B2 => 
                           n20736, ZN => n23998);
   U16203 : OAI211_X1 port map( C1 => n24124, C2 => n24000, A => n23999, B => 
                           n23998, ZN => n5419);
   U16204 : MUX2_X1 port map( A => n21455, B => N241, S => n23184, Z => n5639);
   U16205 : INV_X1 port map( A => N241, ZN => n24098);
   U16206 : OAI222_X1 port map( A1 => n5734, A2 => n22997, B1 => n24098, B2 => 
                           n22996, C1 => n22794, C2 => n22991, ZN => n5644);
   U16207 : INV_X1 port map( A => ADD_WR(0), ZN => n25405);
   U16208 : INV_X1 port map( A => ADD_WR(1), ZN => n25404);
   U16209 : NAND2_X1 port map( A1 => n25405, A2 => n25404, ZN => n24209);
   U16210 : INV_X1 port map( A => n24209, ZN => n24001);
   U16211 : INV_X1 port map( A => ADD_WR(2), ZN => n24202);
   U16212 : INV_X1 port map( A => ADD_WR(3), ZN => n24084);
   U16213 : OAI21_X1 port map( B1 => n24001, B2 => n24202, A => n24084, ZN => 
                           n24130);
   U16214 : AOI22_X1 port map( A1 => n23013, A2 => n21455, B1 => n23029, B2 => 
                           i_31_port, ZN => n24004);
   U16215 : OAI221_X1 port map( B1 => n22779, B2 => n22794, C1 => n967, C2 => 
                           n23007, A => n24004, ZN => U3_U7_Z_31);
   U16216 : NAND2_X1 port map( A1 => n24006, A2 => n24005, ZN => n24085);
   U16217 : NOR2_X1 port map( A1 => n24098, A2 => n23000, ZN => U3_U2_Z_31);
   U16218 : NOR2_X1 port map( A1 => n24099, A2 => n23000, ZN => U3_U2_Z_30);
   U16219 : NOR2_X1 port map( A1 => n24100, A2 => n23000, ZN => U3_U2_Z_29);
   U16220 : NOR2_X1 port map( A1 => n24101, A2 => n23000, ZN => U3_U2_Z_28);
   U16221 : NOR2_X1 port map( A1 => n24102, A2 => n23000, ZN => U3_U2_Z_27);
   U16222 : NOR2_X1 port map( A1 => n24103, A2 => n23000, ZN => U3_U2_Z_26);
   U16223 : NOR2_X1 port map( A1 => n24104, A2 => n23000, ZN => U3_U2_Z_25);
   U16224 : NOR2_X1 port map( A1 => n24105, A2 => n23000, ZN => U3_U2_Z_24);
   U16225 : NOR2_X1 port map( A1 => n24106, A2 => n23000, ZN => U3_U2_Z_23);
   U16226 : NOR2_X1 port map( A1 => n24107, A2 => n23000, ZN => U3_U2_Z_22);
   U16227 : NOR2_X1 port map( A1 => n24108, A2 => n23000, ZN => U3_U2_Z_21);
   U16228 : NOR2_X1 port map( A1 => n24109, A2 => n23000, ZN => U3_U2_Z_20);
   U16229 : NOR2_X1 port map( A1 => n22500, A2 => n23001, ZN => U3_U2_Z_19);
   U16230 : NOR2_X1 port map( A1 => n24111, A2 => n23001, ZN => U3_U2_Z_18);
   U16231 : NOR2_X1 port map( A1 => n24112, A2 => n23001, ZN => U3_U2_Z_17);
   U16232 : INV_X1 port map( A => N226, ZN => n24113);
   U16233 : NOR2_X1 port map( A1 => n24113, A2 => n23001, ZN => U3_U2_Z_16);
   U16234 : NOR2_X1 port map( A1 => n24114, A2 => n23001, ZN => U3_U2_Z_15);
   U16235 : NOR2_X1 port map( A1 => n24115, A2 => n23001, ZN => U3_U2_Z_14);
   U16236 : NOR2_X1 port map( A1 => n24116, A2 => n23001, ZN => U3_U2_Z_13);
   U16237 : NOR2_X1 port map( A1 => n24117, A2 => n23001, ZN => U3_U2_Z_12);
   U16238 : NOR2_X1 port map( A1 => n24118, A2 => n23001, ZN => U3_U2_Z_11);
   U16239 : NOR2_X1 port map( A1 => n22504, A2 => n23001, ZN => U3_U2_Z_10);
   U16240 : NOR2_X1 port map( A1 => n22531, A2 => n23001, ZN => U3_U2_Z_9);
   U16241 : NOR2_X1 port map( A1 => n24121, A2 => n23001, ZN => U3_U2_Z_8);
   U16242 : NOR2_X1 port map( A1 => n24122, A2 => n23002, ZN => U3_U2_Z_7);
   U16243 : NOR2_X1 port map( A1 => n24123, A2 => n23002, ZN => U3_U2_Z_6);
   U16244 : NOR2_X1 port map( A1 => n24124, A2 => n23002, ZN => U3_U2_Z_5);
   U16245 : NAND2_X1 port map( A1 => n24085, A2 => n24138, ZN => n24015);
   U16246 : INV_X1 port map( A => n24015, ZN => n24007);
   U16247 : OAI21_X1 port map( B1 => n24007, B2 => n23004, A => n23034, ZN => 
                           U3_U2_Z_4);
   U16248 : INV_X1 port map( A => ADD_RD1(3), ZN => n24350);
   U16249 : NAND3_X1 port map( A1 => n24008, A2 => n23037, A3 => n22700, ZN => 
                           n24129);
   U16250 : INV_X1 port map( A => n24129, ZN => n24307);
   U16251 : NAND2_X1 port map( A1 => RD1, A2 => n24307, ZN => n24343);
   U16252 : OAI221_X1 port map( B1 => n24290, B2 => n23002, C1 => n24350, C2 =>
                           n24343, A => n23037, ZN => U3_U2_Z_3);
   U16253 : OAI22_X1 port map( A1 => n22796, A2 => n23002, B1 => n24369, B2 => 
                           n24343, ZN => U3_U2_Z_2);
   U16254 : NAND2_X1 port map( A1 => n24085, A2 => n22497, ZN => n24012);
   U16255 : INV_X1 port map( A => n24012, ZN => n24009);
   U16256 : INV_X1 port map( A => ADD_RD1(1), ZN => n24355);
   U16257 : OAI22_X1 port map( A1 => n24009, A2 => n23003, B1 => n24355, B2 => 
                           n24343, ZN => U3_U2_Z_1);
   U16258 : INV_X1 port map( A => ADD_RD1(0), ZN => n24368);
   U16259 : OAI22_X1 port map( A1 => n22505, A2 => n23002, B1 => n24368, B2 => 
                           n24343, ZN => U3_U2_Z_0);
   U16260 : INV_X1 port map( A => N106, ZN => n24096);
   U16261 : OAI22_X1 port map( A1 => n23003, A2 => n22794, B1 => n23034, B2 => 
                           n24096, ZN => U3_U3_Z_31);
   U16262 : INV_X1 port map( A => N105, ZN => n24043);
   U16263 : OAI22_X1 port map( A1 => n23004, A2 => n24045, B1 => n23034, B2 => 
                           n24043, ZN => U3_U3_Z_30);
   U16264 : INV_X1 port map( A => N104, ZN => n24042);
   U16265 : OAI22_X1 port map( A1 => n23003, A2 => n24047, B1 => n24042, B2 => 
                           n23034, ZN => U3_U3_Z_29);
   U16266 : INV_X1 port map( A => N103, ZN => n24041);
   U16267 : OAI22_X1 port map( A1 => n23004, A2 => n22790, B1 => n23034, B2 => 
                           n24041, ZN => U3_U3_Z_28);
   U16268 : INV_X1 port map( A => N102, ZN => n24040);
   U16269 : OAI22_X1 port map( A1 => n23003, A2 => n22789, B1 => n24040, B2 => 
                           n23034, ZN => U3_U3_Z_27);
   U16270 : INV_X1 port map( A => N101, ZN => n24039);
   U16271 : OAI22_X1 port map( A1 => n23004, A2 => n22785, B1 => n23034, B2 => 
                           n24039, ZN => U3_U3_Z_26);
   U16272 : INV_X1 port map( A => N100, ZN => n24038);
   U16273 : OAI22_X1 port map( A1 => n23004, A2 => n22783, B1 => n23034, B2 => 
                           n24038, ZN => U3_U3_Z_25);
   U16274 : INV_X1 port map( A => N99, ZN => n24037);
   U16275 : OAI22_X1 port map( A1 => n23004, A2 => n22981, B1 => n23035, B2 => 
                           n24037, ZN => U3_U3_Z_24);
   U16276 : INV_X1 port map( A => N98, ZN => n24036);
   U16277 : OAI22_X1 port map( A1 => n23004, A2 => n22795, B1 => n23035, B2 => 
                           n24036, ZN => U3_U3_Z_23);
   U16278 : INV_X1 port map( A => N97, ZN => n24035);
   U16279 : OAI22_X1 port map( A1 => n23004, A2 => n22793, B1 => n23035, B2 => 
                           n24035, ZN => U3_U3_Z_22);
   U16280 : INV_X1 port map( A => N96, ZN => n24034);
   U16281 : OAI22_X1 port map( A1 => n23004, A2 => n22786, B1 => n23035, B2 => 
                           n24034, ZN => U3_U3_Z_21);
   U16282 : INV_X1 port map( A => N95, ZN => n24033);
   U16283 : OAI22_X1 port map( A1 => n23004, A2 => n22509, B1 => n23035, B2 => 
                           n24033, ZN => U3_U3_Z_20);
   U16284 : INV_X1 port map( A => N94, ZN => n24032);
   U16285 : OAI22_X1 port map( A1 => n23004, A2 => n24058, B1 => n23035, B2 => 
                           n24032, ZN => U3_U3_Z_19);
   U16286 : INV_X1 port map( A => N93, ZN => n24031);
   U16287 : OAI22_X1 port map( A1 => n23004, A2 => n24060, B1 => n23034, B2 => 
                           n24031, ZN => U3_U3_Z_18);
   U16288 : INV_X1 port map( A => N92, ZN => n24030);
   U16289 : OAI22_X1 port map( A1 => n23004, A2 => n24062, B1 => n23035, B2 => 
                           n24030, ZN => U3_U3_Z_17);
   U16290 : INV_X1 port map( A => N91, ZN => n24029);
   U16291 : OAI22_X1 port map( A1 => n23004, A2 => n22780, B1 => n23035, B2 => 
                           n24029, ZN => U3_U3_Z_16);
   U16292 : INV_X1 port map( A => N90, ZN => n24028);
   U16293 : OAI22_X1 port map( A1 => n23004, A2 => n24065, B1 => n23035, B2 => 
                           n24028, ZN => U3_U3_Z_15);
   U16294 : INV_X1 port map( A => N89, ZN => n24027);
   U16295 : OAI22_X1 port map( A1 => n23003, A2 => n22782, B1 => n23035, B2 => 
                           n24027, ZN => U3_U3_Z_14);
   U16296 : INV_X1 port map( A => N88, ZN => n24026);
   U16297 : OAI22_X1 port map( A1 => n23003, A2 => n22781, B1 => n24026, B2 => 
                           n23035, ZN => U3_U3_Z_13);
   U16298 : INV_X1 port map( A => N87, ZN => n24025);
   U16299 : OAI22_X1 port map( A1 => n23003, A2 => n24069, B1 => n23036, B2 => 
                           n24025, ZN => U3_U3_Z_12);
   U16300 : INV_X1 port map( A => N86, ZN => n24024);
   U16301 : OAI22_X1 port map( A1 => n23003, A2 => n24071, B1 => n24024, B2 => 
                           n23036, ZN => U3_U3_Z_11);
   U16302 : INV_X1 port map( A => N85, ZN => n24023);
   U16303 : OAI22_X1 port map( A1 => n23003, A2 => n24073, B1 => n24023, B2 => 
                           n23036, ZN => U3_U3_Z_10);
   U16304 : INV_X1 port map( A => N84, ZN => n24022);
   U16305 : OAI22_X1 port map( A1 => n23003, A2 => n22539, B1 => n23036, B2 => 
                           n24022, ZN => U3_U3_Z_9);
   U16306 : INV_X1 port map( A => N83, ZN => n24021);
   U16307 : OAI22_X1 port map( A1 => n23004, A2 => n22792, B1 => n23036, B2 => 
                           n24021, ZN => U3_U3_Z_8);
   U16308 : INV_X1 port map( A => N82, ZN => n24020);
   U16309 : OAI22_X1 port map( A1 => n23003, A2 => n22540, B1 => n23036, B2 => 
                           n24020, ZN => U3_U3_Z_7);
   U16310 : INV_X1 port map( A => N81, ZN => n24019);
   U16311 : OAI22_X1 port map( A1 => n23003, A2 => n22791, B1 => n24019, B2 => 
                           n23036, ZN => U3_U3_Z_6);
   U16312 : INV_X1 port map( A => N80, ZN => n24018);
   U16313 : OAI22_X1 port map( A1 => n23003, A2 => n22541, B1 => n23036, B2 => 
                           n24018, ZN => U3_U3_Z_5);
   U16314 : OAI22_X1 port map( A1 => n23003, A2 => n22787, B1 => n23036, B2 => 
                           n24179, ZN => U3_U3_Z_4);
   U16315 : INV_X1 port map( A => N78, ZN => n24292);
   U16316 : OAI22_X1 port map( A1 => n23003, A2 => n22784, B1 => n23035, B2 => 
                           n24292, ZN => U3_U3_Z_3);
   U16317 : INV_X1 port map( A => N77, ZN => n24176);
   U16318 : OAI221_X1 port map( B1 => n23003, B2 => n22983, C1 => n23037, C2 =>
                           n24176, A => n24343, ZN => U3_U3_Z_2);
   U16319 : INV_X1 port map( A => N76, ZN => n24175);
   U16320 : OAI22_X1 port map( A1 => n23003, A2 => n22982, B1 => n23034, B2 => 
                           n24175, ZN => U3_U3_Z_1);
   U16321 : INV_X1 port map( A => N75, ZN => n24125);
   U16322 : OAI221_X1 port map( B1 => n23004, B2 => n22788, C1 => n23037, C2 =>
                           n24125, A => n24343, ZN => U3_U3_Z_0);
   U16323 : NAND2_X1 port map( A1 => n24010, A2 => n23283, ZN => n24011);
   U16324 : OR3_X1 port map( A1 => n23037, A2 => n24011, A3 => N139, ZN => 
                           n24097);
   U16325 : INV_X1 port map( A => n24011, ZN => n24094);
   U16326 : NAND3_X1 port map( A1 => n23016, A2 => n23037, A3 => n24085, ZN => 
                           n24095);
   U16327 : OAI222_X1 port map( A1 => n24125, A2 => n23023, B1 => n22505, B2 =>
                           n23019, C1 => n3046, C2 => n23016, ZN => n5418);
   U16328 : OAI222_X1 port map( A1 => n24176, A2 => n23023, B1 => n22797, B2 =>
                           n23019, C1 => n3045, C2 => n23018, ZN => n5417);
   U16329 : NAND2_X1 port map( A1 => n24012, A2 => n23037, ZN => n24013);
   U16330 : MUX2_X1 port map( A => n3044, B => n24013, S => n23016, Z => n24014
                           );
   U16331 : OAI21_X1 port map( B1 => n24175, B2 => n23025, A => n24014, ZN => 
                           n5416);
   U16332 : OAI222_X1 port map( A1 => n24292, A2 => n23023, B1 => n24290, B2 =>
                           n23019, C1 => n3043, C2 => n23018, ZN => n5415);
   U16333 : NAND2_X1 port map( A1 => n24015, A2 => n23036, ZN => n24016);
   U16334 : MUX2_X1 port map( A => n994, B => n24016, S => n23016, Z => n24017)
                           ;
   U16335 : OAI21_X1 port map( B1 => n24179, B2 => n23025, A => n24017, ZN => 
                           n3366);
   U16336 : OAI222_X1 port map( A1 => n23025, A2 => n24018, B1 => n24124, B2 =>
                           n23019, C1 => n993, C2 => n23018, ZN => n3365);
   U16337 : OAI222_X1 port map( A1 => n23025, A2 => n24019, B1 => n24123, B2 =>
                           n23019, C1 => n992, C2 => n23018, ZN => n3364);
   U16338 : OAI222_X1 port map( A1 => n23025, A2 => n24020, B1 => n24122, B2 =>
                           n23019, C1 => n991, C2 => n23018, ZN => n3363);
   U16339 : OAI222_X1 port map( A1 => n23025, A2 => n24021, B1 => n24121, B2 =>
                           n23019, C1 => n990, C2 => n23018, ZN => n3362);
   U16340 : OAI222_X1 port map( A1 => n23025, A2 => n24022, B1 => n22531, B2 =>
                           n23019, C1 => n989, C2 => n23018, ZN => n3361);
   U16341 : OAI222_X1 port map( A1 => n23024, A2 => n24025, B1 => n24117, B2 =>
                           n23019, C1 => n986, C2 => n23017, ZN => n3358);
   U16342 : OAI222_X1 port map( A1 => n23024, A2 => n24027, B1 => n24115, B2 =>
                           n23020, C1 => n984, C2 => n23017, ZN => n3356);
   U16343 : OAI222_X1 port map( A1 => n23024, A2 => n24028, B1 => n24114, B2 =>
                           n23020, C1 => n983, C2 => n23017, ZN => n3355);
   U16344 : OAI222_X1 port map( A1 => n23024, A2 => n24029, B1 => n24113, B2 =>
                           n23020, C1 => n982, C2 => n23017, ZN => n3354);
   U16345 : OAI222_X1 port map( A1 => n23024, A2 => n24030, B1 => n24112, B2 =>
                           n23020, C1 => n981, C2 => n23017, ZN => n3353);
   U16346 : OAI222_X1 port map( A1 => n23024, A2 => n24031, B1 => n24111, B2 =>
                           n23020, C1 => n980, C2 => n23017, ZN => n3352);
   U16347 : OAI222_X1 port map( A1 => n23024, A2 => n24032, B1 => n22500, B2 =>
                           n23020, C1 => n979, C2 => n23017, ZN => n3351);
   U16348 : OAI222_X1 port map( A1 => n23024, A2 => n24033, B1 => n24109, B2 =>
                           n23020, C1 => n978, C2 => n23017, ZN => n3350);
   U16349 : OAI222_X1 port map( A1 => n23024, A2 => n24034, B1 => n24108, B2 =>
                           n23020, C1 => n977, C2 => n23017, ZN => n3349);
   U16350 : OAI222_X1 port map( A1 => n23023, A2 => n24035, B1 => n24107, B2 =>
                           n23020, C1 => n976, C2 => n23016, ZN => n3348);
   U16351 : OAI222_X1 port map( A1 => n23023, A2 => n24036, B1 => n24106, B2 =>
                           n23020, C1 => n975, C2 => n23016, ZN => n3347);
   U16352 : OAI222_X1 port map( A1 => n23023, A2 => n24037, B1 => n24105, B2 =>
                           n23020, C1 => n974, C2 => n23016, ZN => n3346);
   U16353 : OAI222_X1 port map( A1 => n23023, A2 => n24038, B1 => n24104, B2 =>
                           n23020, C1 => n973, C2 => n23016, ZN => n3345);
   U16354 : OAI222_X1 port map( A1 => n23023, A2 => n24039, B1 => n24103, B2 =>
                           n23021, C1 => n972, C2 => n23016, ZN => n3344);
   U16355 : OAI222_X1 port map( A1 => n23023, A2 => n24040, B1 => n24102, B2 =>
                           n23021, C1 => n971, C2 => n23016, ZN => n3343);
   U16356 : OAI222_X1 port map( A1 => n23023, A2 => n24042, B1 => n24100, B2 =>
                           n23021, C1 => n969, C2 => n23016, ZN => n3341);
   U16357 : OAI222_X1 port map( A1 => n23023, A2 => n24043, B1 => n24099, B2 =>
                           n23021, C1 => n968, C2 => n23016, ZN => n3340);
   U16358 : AOI22_X1 port map( A1 => n23011, A2 => n21453, B1 => n23029, B2 => 
                           i_30_port, ZN => n24044);
   U16359 : OAI221_X1 port map( B1 => n22777, B2 => n24045, C1 => n968, C2 => 
                           n23007, A => n24044, ZN => U3_U7_Z_30);
   U16360 : AOI22_X1 port map( A1 => n23013, A2 => n21449, B1 => n23029, B2 => 
                           i_29_port, ZN => n24046);
   U16361 : OAI221_X1 port map( B1 => n22778, B2 => n24047, C1 => n969, C2 => 
                           n23007, A => n24046, ZN => U3_U7_Z_29);
   U16362 : AOI22_X1 port map( A1 => n23011, A2 => n21446, B1 => n23028, B2 => 
                           i_28_port, ZN => n24048);
   U16363 : OAI221_X1 port map( B1 => n22779, B2 => n22790, C1 => n970, C2 => 
                           n23007, A => n24048, ZN => U3_U7_Z_28);
   U16364 : AOI22_X1 port map( A1 => n22769, A2 => n21442, B1 => n23029, B2 => 
                           i_27_port, ZN => n24049);
   U16365 : OAI221_X1 port map( B1 => n22777, B2 => n22789, C1 => n971, C2 => 
                           n23007, A => n24049, ZN => U3_U7_Z_27);
   U16366 : AOI22_X1 port map( A1 => n23013, A2 => n21441, B1 => n23028, B2 => 
                           i_26_port, ZN => n24050);
   U16367 : OAI221_X1 port map( B1 => n22779, B2 => n22785, C1 => n972, C2 => 
                           n23007, A => n24050, ZN => U3_U7_Z_26);
   U16368 : AOI22_X1 port map( A1 => n23011, A2 => n21439, B1 => n23029, B2 => 
                           i_25_port, ZN => n24051);
   U16369 : OAI221_X1 port map( B1 => n22779, B2 => n22783, C1 => n973, C2 => 
                           n23007, A => n24051, ZN => U3_U7_Z_25);
   U16370 : AOI22_X1 port map( A1 => n22769, A2 => n21437, B1 => n23028, B2 => 
                           i_24_port, ZN => n24052);
   U16371 : OAI221_X1 port map( B1 => n22779, B2 => n22981, C1 => n974, C2 => 
                           n23007, A => n24052, ZN => U3_U7_Z_24);
   U16372 : AOI22_X1 port map( A1 => n23013, A2 => n21434, B1 => n23028, B2 => 
                           i_23_port, ZN => n24053);
   U16373 : AOI22_X1 port map( A1 => n23011, A2 => n21433, B1 => n23028, B2 => 
                           i_22_port, ZN => n24054);
   U16374 : AOI22_X1 port map( A1 => n23013, A2 => n21436, B1 => n23028, B2 => 
                           i_21_port, ZN => n24055);
   U16375 : OAI221_X1 port map( B1 => n22779, B2 => n22786, C1 => n977, C2 => 
                           n23007, A => n24055, ZN => U3_U7_Z_21);
   U16376 : AOI22_X1 port map( A1 => n23011, A2 => n21435, B1 => n23029, B2 => 
                           i_20_port, ZN => n24056);
   U16377 : OAI221_X1 port map( B1 => n22778, B2 => n22509, C1 => n978, C2 => 
                           n23007, A => n24056, ZN => U3_U7_Z_20);
   U16378 : AOI22_X1 port map( A1 => n23013, A2 => n21030, B1 => n23028, B2 => 
                           i_19_port, ZN => n24057);
   U16379 : OAI221_X1 port map( B1 => n22770, B2 => n24058, C1 => n979, C2 => 
                           n23008, A => n24057, ZN => U3_U7_Z_19);
   U16380 : AOI22_X1 port map( A1 => n23013, A2 => n21430, B1 => n23029, B2 => 
                           i_18_port, ZN => n24059);
   U16381 : AOI22_X1 port map( A1 => n23011, A2 => n21431, B1 => n23029, B2 => 
                           i_17_port, ZN => n24061);
   U16382 : OAI221_X1 port map( B1 => n22770, B2 => n24062, C1 => n981, C2 => 
                           n23008, A => n24061, ZN => U3_U7_Z_17);
   U16383 : AOI22_X1 port map( A1 => n22769, A2 => n21432, B1 => n23028, B2 => 
                           i_16_port, ZN => n24063);
   U16384 : OAI221_X1 port map( B1 => n22770, B2 => n22780, C1 => n982, C2 => 
                           n23008, A => n24063, ZN => U3_U7_Z_16);
   U16385 : AOI22_X1 port map( A1 => n23011, A2 => n21428, B1 => n23028, B2 => 
                           i_15_port, ZN => n24064);
   U16386 : OAI221_X1 port map( B1 => n22771, B2 => n24065, C1 => n983, C2 => 
                           n23008, A => n24064, ZN => U3_U7_Z_15);
   U16387 : AOI22_X1 port map( A1 => n23013, A2 => n21029, B1 => n23029, B2 => 
                           i_14_port, ZN => n24066);
   U16388 : OAI221_X1 port map( B1 => n22773, B2 => n22782, C1 => n984, C2 => 
                           n23008, A => n24066, ZN => U3_U7_Z_14);
   U16389 : AOI22_X1 port map( A1 => n23013, A2 => n21426, B1 => n23028, B2 => 
                           i_13_port, ZN => n24067);
   U16390 : OAI221_X1 port map( B1 => n22774, B2 => n22781, C1 => n985, C2 => 
                           n23008, A => n24067, ZN => U3_U7_Z_13);
   U16391 : AOI22_X1 port map( A1 => n22769, A2 => n21427, B1 => n23029, B2 => 
                           i_12_port, ZN => n24068);
   U16392 : OAI221_X1 port map( B1 => n22773, B2 => n24069, C1 => n986, C2 => 
                           n23008, A => n24068, ZN => U3_U7_Z_12);
   U16393 : AOI22_X1 port map( A1 => n23011, A2 => n21028, B1 => n23028, B2 => 
                           i_11_port, ZN => n24070);
   U16394 : OAI221_X1 port map( B1 => n22773, B2 => n24071, C1 => n987, C2 => 
                           n23008, A => n24070, ZN => U3_U7_Z_11);
   U16395 : AOI22_X1 port map( A1 => n23013, A2 => n21425, B1 => n23028, B2 => 
                           i_10_port, ZN => n24072);
   U16396 : OAI221_X1 port map( B1 => n22773, B2 => n24073, C1 => n988, C2 => 
                           n23008, A => n24072, ZN => U3_U7_Z_10);
   U16397 : AOI22_X1 port map( A1 => n23013, A2 => n21027, B1 => n23028, B2 => 
                           i_9_port, ZN => n24074);
   U16398 : OAI221_X1 port map( B1 => n22774, B2 => n22539, C1 => n989, C2 => 
                           n23008, A => n24074, ZN => U3_U7_Z_9);
   U16399 : AOI22_X1 port map( A1 => n23012, A2 => n21424, B1 => n23029, B2 => 
                           i_8_port, ZN => n24075);
   U16400 : OAI221_X1 port map( B1 => n22775, B2 => n22792, C1 => n990, C2 => 
                           n23008, A => n24075, ZN => U3_U7_Z_8);
   U16401 : AOI22_X1 port map( A1 => n23012, A2 => n21423, B1 => n23027, B2 => 
                           i_7_port, ZN => n24076);
   U16402 : OAI221_X1 port map( B1 => n23015, B2 => n22540, C1 => n991, C2 => 
                           n23009, A => n24076, ZN => U3_U7_Z_7);
   U16403 : AOI22_X1 port map( A1 => n23012, A2 => n21421, B1 => n23027, B2 => 
                           i_6_port, ZN => n24077);
   U16404 : OAI221_X1 port map( B1 => n23015, B2 => n22791, C1 => n992, C2 => 
                           n23009, A => n24077, ZN => U3_U7_Z_6);
   U16405 : AOI22_X1 port map( A1 => n23012, A2 => n21422, B1 => n23027, B2 => 
                           i_5_port, ZN => n24078);
   U16406 : OAI221_X1 port map( B1 => n23015, B2 => n22541, C1 => n993, C2 => 
                           n23009, A => n24078, ZN => U3_U7_Z_5);
   U16407 : AOI22_X1 port map( A1 => n23012, A2 => n21420, B1 => n23027, B2 => 
                           i_4_port, ZN => n24079);
   U16408 : OAI221_X1 port map( B1 => n23015, B2 => n22787, C1 => n994, C2 => 
                           n23009, A => n24079, ZN => U3_U7_Z_4);
   U16409 : AOI22_X1 port map( A1 => n23014, A2 => n21418, B1 => n23030, B2 => 
                           i_3_port, ZN => n24080);
   U16410 : AOI22_X1 port map( A1 => n23014, A2 => n21419, B1 => n23030, B2 => 
                           n24143, ZN => n24081);
   U16411 : OAI221_X1 port map( B1 => n24090, B2 => n22983, C1 => n3045, C2 => 
                           n23009, A => n24081, ZN => U3_U7_Z_2);
   U16412 : AOI22_X1 port map( A1 => n22489, A2 => n21417, B1 => n22502, B2 => 
                           i_1_port, ZN => n24082);
   U16413 : OAI221_X1 port map( B1 => n24090, B2 => n22982, C1 => n3044, C2 => 
                           n23009, A => n24082, ZN => U3_U7_Z_1);
   U16414 : AOI22_X1 port map( A1 => n22489, A2 => n21416, B1 => n22502, B2 => 
                           i_0_port, ZN => n24083);
   U16415 : OAI221_X1 port map( B1 => n24090, B2 => n22788, C1 => n3046, C2 => 
                           n23009, A => n24083, ZN => U3_U7_Z_0);
   U16416 : NOR2_X1 port map( A1 => n22546, A2 => n24084, ZN => U3_U8_Z_3);
   U16417 : NAND2_X1 port map( A1 => n24085, A2 => SIGRETURN, ZN => n24091);
   U16418 : NOR2_X1 port map( A1 => n5700, A2 => n24086, ZN => n24088);
   U16419 : AOI211_X1 port map( C1 => n22510, C2 => n24088, A => n22489, B => 
                           n22502, ZN => n24089);
   U16420 : OAI211_X1 port map( C1 => n24202, C2 => n22545, A => n24091, B => 
                           n24089, ZN => U3_U8_Z_2);
   U16421 : OAI211_X1 port map( C1 => n25404, C2 => n22546, A => n22507, B => 
                           n24092, ZN => n20764);
   U16422 : OAI21_X1 port map( B1 => n25405, B2 => n22545, A => n24093, ZN => 
                           U3_U8_Z_0);
   U16423 : OAI222_X1 port map( A1 => n23024, A2 => n24096, B1 => n24098, B2 =>
                           n23021, C1 => n967, C2 => n23017, ZN => n3339);
   U16424 : NOR2_X1 port map( A1 => n23031, A2 => n24098, ZN => U3_U1_Z_31);
   U16425 : NOR2_X1 port map( A1 => n23031, A2 => n24099, ZN => U3_U1_Z_30);
   U16426 : NOR2_X1 port map( A1 => n23031, A2 => n24100, ZN => U3_U1_Z_29);
   U16427 : NOR2_X1 port map( A1 => n23031, A2 => n24101, ZN => U3_U1_Z_28);
   U16428 : NOR2_X1 port map( A1 => n23031, A2 => n24102, ZN => U3_U1_Z_27);
   U16429 : NOR2_X1 port map( A1 => n23031, A2 => n24103, ZN => U3_U1_Z_26);
   U16430 : NOR2_X1 port map( A1 => n23031, A2 => n24104, ZN => U3_U1_Z_25);
   U16431 : NOR2_X1 port map( A1 => n23031, A2 => n24105, ZN => U3_U1_Z_24);
   U16432 : NOR2_X1 port map( A1 => n24107, A2 => n23031, ZN => U3_U1_Z_22);
   U16433 : NOR2_X1 port map( A1 => n23031, A2 => n24108, ZN => U3_U1_Z_21);
   U16434 : NOR2_X1 port map( A1 => n23031, A2 => n24109, ZN => U3_U1_Z_20);
   U16435 : NOR2_X1 port map( A1 => n23031, A2 => n24110, ZN => U3_U1_Z_19);
   U16436 : NOR2_X1 port map( A1 => n23031, A2 => n24111, ZN => U3_U1_Z_18);
   U16437 : NOR2_X1 port map( A1 => n23031, A2 => n24112, ZN => U3_U1_Z_17);
   U16438 : NOR2_X1 port map( A1 => n23031, A2 => n24113, ZN => U3_U1_Z_16);
   U16439 : NOR2_X1 port map( A1 => n23031, A2 => n24116, ZN => U3_U1_Z_13);
   U16440 : NOR2_X1 port map( A1 => n23031, A2 => n24117, ZN => U3_U1_Z_12);
   U16441 : NOR2_X1 port map( A1 => n23031, A2 => n24119, ZN => U3_U1_Z_10);
   U16442 : NOR2_X1 port map( A1 => n23031, A2 => n24120, ZN => U3_U1_Z_9);
   U16443 : NOR2_X1 port map( A1 => n23031, A2 => n24121, ZN => U3_U1_Z_8);
   U16444 : NOR2_X1 port map( A1 => n23031, A2 => n24138, ZN => U3_U1_Z_4);
   U16445 : OAI21_X1 port map( B1 => n23031, B2 => n24183, A => n23034, ZN => 
                           U3_U1_Z_2);
   U16446 : OAI21_X1 port map( B1 => n23031, B2 => n24184, A => n23034, ZN => 
                           U3_U1_Z_1);
   U16447 : NOR2_X1 port map( A1 => n23031, A2 => n24185, ZN => U3_U1_Z_0);
   U16448 : INV_X1 port map( A => n16601, ZN => n24286);
   U16449 : NAND2_X1 port map( A1 => n22490, A2 => n24175, ZN => n24297);
   U16450 : NAND3_X1 port map( A1 => n22689, A2 => n24179, A3 => n24292, ZN => 
                           n24203);
   U16451 : NAND3_X1 port map( A1 => n22532, A2 => n22497, A3 => n22505, ZN => 
                           n24296);
   U16452 : INV_X1 port map( A => n22545, ZN => n24128);
   U16453 : NAND3_X1 port map( A1 => n22695, A2 => n24138, A3 => n24290, ZN => 
                           n24198);
   U16454 : NOR2_X1 port map( A1 => n24202, A2 => n24129, ZN => n24132);
   U16455 : INV_X1 port map( A => n24130, ZN => n24131);
   U16456 : AOI21_X1 port map( B1 => n24132, B2 => n22485, A => RESET, ZN => 
                           n24133);
   U16457 : OAI221_X1 port map( B1 => n24297, B2 => n24203, C1 => n24296, C2 =>
                           n24198, A => n24133, ZN => n24134);
   U16458 : INV_X1 port map( A => n24134, ZN => n24135);
   U16459 : MUX2_X1 port map( A => n24286, B => n22229, S => n23056, Z => n5158
                           );
   U16460 : INV_X1 port map( A => n16602, ZN => n24272);
   U16461 : MUX2_X1 port map( A => n24272, B => n22230, S => n23056, Z => n5157
                           );
   U16462 : INV_X1 port map( A => n16603, ZN => n24270);
   U16463 : MUX2_X1 port map( A => n24270, B => n22231, S => n23056, Z => n5156
                           );
   U16464 : INV_X1 port map( A => n16604, ZN => n24268);
   U16465 : MUX2_X1 port map( A => n24268, B => n22232, S => n23056, Z => n5155
                           );
   U16466 : INV_X1 port map( A => n16605, ZN => n24266);
   U16467 : MUX2_X1 port map( A => n24266, B => n22233, S => n23056, Z => n5154
                           );
   U16468 : INV_X1 port map( A => n16606, ZN => n24264);
   U16469 : MUX2_X1 port map( A => n24264, B => n22234, S => n23056, Z => n5153
                           );
   U16470 : INV_X1 port map( A => n16607, ZN => n24262);
   U16471 : MUX2_X1 port map( A => n24262, B => n22227, S => n23056, Z => n5152
                           );
   U16472 : INV_X1 port map( A => n16608, ZN => n24260);
   U16473 : MUX2_X1 port map( A => n24260, B => n22235, S => n23056, Z => n5151
                           );
   U16474 : INV_X1 port map( A => n16609, ZN => n24258);
   U16475 : MUX2_X1 port map( A => n24258, B => n22236, S => n23056, Z => n5150
                           );
   U16476 : INV_X1 port map( A => n16610, ZN => n24256);
   U16477 : MUX2_X1 port map( A => n24256, B => n22237, S => n23056, Z => n5149
                           );
   U16478 : INV_X1 port map( A => n16611, ZN => n24254);
   U16479 : MUX2_X1 port map( A => n24254, B => n22238, S => n23056, Z => n5148
                           );
   U16480 : INV_X1 port map( A => n16612, ZN => n24252);
   U16481 : MUX2_X1 port map( A => n24252, B => n22239, S => n23056, Z => n5147
                           );
   U16482 : INV_X1 port map( A => n16613, ZN => n24250);
   U16483 : MUX2_X1 port map( A => n24250, B => n22240, S => n23057, Z => n5146
                           );
   U16484 : INV_X1 port map( A => n16614, ZN => n24248);
   U16485 : MUX2_X1 port map( A => n24248, B => n22241, S => n23057, Z => n5145
                           );
   U16486 : INV_X1 port map( A => n16615, ZN => n24246);
   U16487 : MUX2_X1 port map( A => n24246, B => n22242, S => n23057, Z => n5144
                           );
   U16488 : INV_X1 port map( A => n16616, ZN => n24244);
   U16489 : MUX2_X1 port map( A => n24244, B => n22243, S => n23057, Z => n5143
                           );
   U16490 : INV_X1 port map( A => n16617, ZN => n24242);
   U16491 : MUX2_X1 port map( A => n24242, B => n22244, S => n23057, Z => n5142
                           );
   U16492 : INV_X1 port map( A => n16618, ZN => n24240);
   U16493 : MUX2_X1 port map( A => n24240, B => n22245, S => n23057, Z => n5141
                           );
   U16494 : INV_X1 port map( A => n16619, ZN => n24238);
   U16495 : MUX2_X1 port map( A => n24238, B => n22228, S => n23057, Z => n5140
                           );
   U16496 : INV_X1 port map( A => n16620, ZN => n24236);
   U16497 : MUX2_X1 port map( A => n24236, B => n22246, S => n23057, Z => n5139
                           );
   U16498 : INV_X1 port map( A => n16621, ZN => n24234);
   U16499 : MUX2_X1 port map( A => n24234, B => n22247, S => n23057, Z => n5138
                           );
   U16500 : INV_X1 port map( A => n16622, ZN => n24232);
   U16501 : MUX2_X1 port map( A => n24232, B => n22248, S => n23057, Z => n5137
                           );
   U16502 : INV_X1 port map( A => n16623, ZN => n24230);
   U16503 : MUX2_X1 port map( A => n24230, B => n22249, S => n23057, Z => n5136
                           );
   U16504 : INV_X1 port map( A => n16624, ZN => n24228);
   U16505 : MUX2_X1 port map( A => n24228, B => n22261, S => n23057, Z => n5135
                           );
   U16506 : INV_X1 port map( A => n16625, ZN => n24226);
   U16507 : MUX2_X1 port map( A => n24226, B => n22250, S => n23058, Z => n5134
                           );
   U16508 : INV_X1 port map( A => n16626, ZN => n24224);
   U16509 : MUX2_X1 port map( A => n24224, B => n22251, S => n23058, Z => n5133
                           );
   U16510 : INV_X1 port map( A => n16627, ZN => n24222);
   U16511 : MUX2_X1 port map( A => n24222, B => n22252, S => n23058, Z => n5132
                           );
   U16512 : INV_X1 port map( A => n16628, ZN => n24220);
   U16513 : MUX2_X1 port map( A => n24220, B => n22253, S => n23058, Z => n5131
                           );
   U16514 : INV_X1 port map( A => n16629, ZN => n24218);
   U16515 : MUX2_X1 port map( A => n24218, B => n22254, S => n23058, Z => n5130
                           );
   U16516 : INV_X1 port map( A => n16630, ZN => n24216);
   U16517 : MUX2_X1 port map( A => n24216, B => n22262, S => n23058, Z => n5129
                           );
   U16518 : INV_X1 port map( A => n16631, ZN => n24214);
   U16519 : MUX2_X1 port map( A => n24214, B => n22255, S => n23058, Z => n5128
                           );
   U16520 : INV_X1 port map( A => n16632, ZN => n24212);
   U16521 : MUX2_X1 port map( A => n24212, B => n22256, S => n23058, Z => n5127
                           );
   U16522 : INV_X1 port map( A => n16633, ZN => n24211);
   U16523 : MUX2_X1 port map( A => n24211, B => n22226, S => n23058, Z => n5126
                           );
   U16524 : INV_X1 port map( A => n16634, ZN => n24213);
   U16525 : MUX2_X1 port map( A => n24213, B => n22257, S => n23058, Z => n5125
                           );
   U16526 : INV_X1 port map( A => n16635, ZN => n24215);
   U16527 : MUX2_X1 port map( A => n24215, B => n22258, S => n23058, Z => n5124
                           );
   U16528 : INV_X1 port map( A => n16636, ZN => n24217);
   U16529 : MUX2_X1 port map( A => n24217, B => n22263, S => n23058, Z => n5123
                           );
   U16530 : INV_X1 port map( A => n16637, ZN => n24219);
   U16531 : MUX2_X1 port map( A => n24219, B => n22264, S => n23059, Z => n5122
                           );
   U16532 : INV_X1 port map( A => n16638, ZN => n24221);
   U16533 : MUX2_X1 port map( A => n24221, B => n22265, S => n23059, Z => n5121
                           );
   U16534 : INV_X1 port map( A => n16639, ZN => n24223);
   U16535 : MUX2_X1 port map( A => n24223, B => n22266, S => n23059, Z => n5120
                           );
   U16536 : INV_X1 port map( A => n16640, ZN => n24225);
   U16537 : MUX2_X1 port map( A => n24225, B => n22267, S => n23059, Z => n5119
                           );
   U16538 : INV_X1 port map( A => n16641, ZN => n24227);
   U16539 : MUX2_X1 port map( A => n24227, B => n22268, S => n23059, Z => n5118
                           );
   U16540 : INV_X1 port map( A => n16642, ZN => n24229);
   U16541 : MUX2_X1 port map( A => n24229, B => n22259, S => n23059, Z => n5117
                           );
   U16542 : INV_X1 port map( A => n16643, ZN => n24231);
   U16543 : MUX2_X1 port map( A => n24231, B => n22269, S => n23059, Z => n5116
                           );
   U16544 : INV_X1 port map( A => n16644, ZN => n24233);
   U16545 : MUX2_X1 port map( A => n24233, B => n22270, S => n23059, Z => n5115
                           );
   U16546 : INV_X1 port map( A => n16645, ZN => n24235);
   U16547 : MUX2_X1 port map( A => n24235, B => n22271, S => n23059, Z => n5114
                           );
   U16548 : INV_X1 port map( A => n16646, ZN => n24237);
   U16549 : MUX2_X1 port map( A => n24237, B => n22272, S => n23059, Z => n5113
                           );
   U16550 : INV_X1 port map( A => n16647, ZN => n24239);
   U16551 : MUX2_X1 port map( A => n24239, B => n22273, S => n23059, Z => n5112
                           );
   U16552 : INV_X1 port map( A => n16648, ZN => n24241);
   U16553 : MUX2_X1 port map( A => n24241, B => n22274, S => n23059, Z => n5111
                           );
   U16554 : INV_X1 port map( A => n16649, ZN => n24243);
   U16555 : MUX2_X1 port map( A => n24243, B => n22275, S => n23060, Z => n5110
                           );
   U16556 : INV_X1 port map( A => n16650, ZN => n24245);
   U16557 : MUX2_X1 port map( A => n24245, B => n22276, S => n23060, Z => n5109
                           );
   U16558 : INV_X1 port map( A => n16651, ZN => n24247);
   U16559 : MUX2_X1 port map( A => n24247, B => n22277, S => n23060, Z => n5108
                           );
   U16560 : INV_X1 port map( A => n16652, ZN => n24249);
   U16561 : MUX2_X1 port map( A => n24249, B => n22278, S => n23060, Z => n5107
                           );
   U16562 : INV_X1 port map( A => n16653, ZN => n24251);
   U16563 : MUX2_X1 port map( A => n24251, B => n22279, S => n23060, Z => n5106
                           );
   U16564 : INV_X1 port map( A => n16654, ZN => n24253);
   U16565 : MUX2_X1 port map( A => n24253, B => n22260, S => n23060, Z => n5105
                           );
   U16566 : INV_X1 port map( A => n16655, ZN => n24255);
   U16567 : MUX2_X1 port map( A => n24255, B => n22280, S => n23060, Z => n5104
                           );
   U16568 : INV_X1 port map( A => n16656, ZN => n24257);
   U16569 : MUX2_X1 port map( A => n24257, B => n22281, S => n23060, Z => n5103
                           );
   U16570 : INV_X1 port map( A => n16657, ZN => n24259);
   U16571 : MUX2_X1 port map( A => n24259, B => n22282, S => n23060, Z => n5102
                           );
   U16572 : INV_X1 port map( A => n16658, ZN => n24261);
   U16573 : MUX2_X1 port map( A => n24261, B => n22283, S => n23060, Z => n5101
                           );
   U16574 : INV_X1 port map( A => n16659, ZN => n24263);
   U16575 : MUX2_X1 port map( A => n24263, B => n22284, S => n23060, Z => n5100
                           );
   U16576 : INV_X1 port map( A => n16660, ZN => n24265);
   U16577 : MUX2_X1 port map( A => n24265, B => n22285, S => n23060, Z => n5099
                           );
   U16578 : INV_X1 port map( A => n16661, ZN => n24267);
   U16579 : MUX2_X1 port map( A => n24267, B => n22286, S => n23061, Z => n5098
                           );
   U16580 : INV_X1 port map( A => n16662, ZN => n24269);
   U16581 : MUX2_X1 port map( A => n24269, B => n22287, S => n23061, Z => n5097
                           );
   U16582 : INV_X1 port map( A => n16663, ZN => n24271);
   U16583 : MUX2_X1 port map( A => n24271, B => n22288, S => n23061, Z => n5096
                           );
   U16584 : INV_X1 port map( A => n16664, ZN => n24273);
   U16585 : MUX2_X1 port map( A => n24273, B => n22289, S => n23061, Z => n5095
                           );
   U16586 : NAND3_X1 port map( A1 => n22532, A2 => n22506, A3 => n22497, ZN => 
                           n24295);
   U16587 : NAND3_X1 port map( A1 => n22694, A2 => n24179, A3 => n24292, ZN => 
                           n24190);
   U16588 : OAI221_X1 port map( B1 => n24295, B2 => n24198, C1 => n24297, C2 =>
                           n24190, A => n23284, ZN => n24136);
   U16589 : INV_X1 port map( A => n24136, ZN => n24137);
   U16590 : MUX2_X1 port map( A => n24286, B => n22057, S => n23064, Z => n5094
                           );
   U16591 : MUX2_X1 port map( A => n24272, B => n22182, S => n23064, Z => n5093
                           );
   U16592 : MUX2_X1 port map( A => n24270, B => n22056, S => n23064, Z => n5092
                           );
   U16593 : MUX2_X1 port map( A => n24268, B => n22179, S => n23064, Z => n5091
                           );
   U16594 : MUX2_X1 port map( A => n24266, B => n22036, S => n23064, Z => n5090
                           );
   U16595 : MUX2_X1 port map( A => n24264, B => n22055, S => n23064, Z => n5089
                           );
   U16596 : MUX2_X1 port map( A => n24262, B => n22175, S => n23064, Z => n5088
                           );
   U16597 : MUX2_X1 port map( A => n24260, B => n22173, S => n23064, Z => n5087
                           );
   U16598 : MUX2_X1 port map( A => n24258, B => n22172, S => n23064, Z => n5086
                           );
   U16599 : MUX2_X1 port map( A => n24256, B => n22170, S => n23064, Z => n5085
                           );
   U16600 : MUX2_X1 port map( A => n24254, B => n22168, S => n23064, Z => n5084
                           );
   U16601 : MUX2_X1 port map( A => n24252, B => n22053, S => n23064, Z => n5083
                           );
   U16602 : MUX2_X1 port map( A => n24250, B => n22165, S => n23065, Z => n5082
                           );
   U16603 : MUX2_X1 port map( A => n24248, B => n22164, S => n23065, Z => n5081
                           );
   U16604 : MUX2_X1 port map( A => n24246, B => n22162, S => n23065, Z => n5080
                           );
   U16605 : MUX2_X1 port map( A => n24244, B => n22051, S => n23065, Z => n5079
                           );
   U16606 : MUX2_X1 port map( A => n24242, B => n22049, S => n23065, Z => n5078
                           );
   U16607 : MUX2_X1 port map( A => n24240, B => n22047, S => n23065, Z => n5077
                           );
   U16608 : MUX2_X1 port map( A => n24238, B => n22045, S => n23065, Z => n5076
                           );
   U16609 : MUX2_X1 port map( A => n24236, B => n22043, S => n23065, Z => n5075
                           );
   U16610 : MUX2_X1 port map( A => n24234, B => n22159, S => n23065, Z => n5074
                           );
   U16611 : MUX2_X1 port map( A => n24232, B => n22158, S => n23065, Z => n5073
                           );
   U16612 : MUX2_X1 port map( A => n24230, B => n22156, S => n23065, Z => n5072
                           );
   U16613 : MUX2_X1 port map( A => n24228, B => n22155, S => n23065, Z => n5071
                           );
   U16614 : MUX2_X1 port map( A => n24226, B => n22040, S => n23066, Z => n5070
                           );
   U16615 : MUX2_X1 port map( A => n24224, B => n22152, S => n23066, Z => n5069
                           );
   U16616 : MUX2_X1 port map( A => n24222, B => n22150, S => n23066, Z => n5068
                           );
   U16617 : MUX2_X1 port map( A => n24220, B => n22039, S => n23066, Z => n5067
                           );
   U16618 : MUX2_X1 port map( A => n24218, B => n22147, S => n23066, Z => n5066
                           );
   U16619 : MUX2_X1 port map( A => n24216, B => n22145, S => n23066, Z => n5065
                           );
   U16620 : MUX2_X1 port map( A => n24214, B => n22038, S => n23066, Z => n5064
                           );
   U16621 : MUX2_X1 port map( A => n24212, B => n22143, S => n23066, Z => n5063
                           );
   U16622 : MUX2_X1 port map( A => n24211, B => n22291, S => n23066, Z => n5062
                           );
   U16623 : MUX2_X1 port map( A => n24213, B => n22037, S => n23066, Z => n5061
                           );
   U16624 : MUX2_X1 port map( A => n24215, B => n22144, S => n23066, Z => n5060
                           );
   U16625 : MUX2_X1 port map( A => n24217, B => n22146, S => n23066, Z => n5059
                           );
   U16626 : MUX2_X1 port map( A => n24219, B => n22148, S => n23067, Z => n5058
                           );
   U16627 : MUX2_X1 port map( A => n24221, B => n22149, S => n23067, Z => n5057
                           );
   U16628 : MUX2_X1 port map( A => n24223, B => n22151, S => n23067, Z => n5056
                           );
   U16629 : MUX2_X1 port map( A => n24225, B => n22153, S => n23067, Z => n5055
                           );
   U16630 : MUX2_X1 port map( A => n24227, B => n22154, S => n23067, Z => n5054
                           );
   U16631 : MUX2_X1 port map( A => n24229, B => n22041, S => n23067, Z => n5053
                           );
   U16632 : MUX2_X1 port map( A => n24231, B => n22157, S => n23067, Z => n5052
                           );
   U16633 : MUX2_X1 port map( A => n24233, B => n22042, S => n23067, Z => n5051
                           );
   U16634 : MUX2_X1 port map( A => n24235, B => n22160, S => n23067, Z => n5050
                           );
   U16635 : MUX2_X1 port map( A => n24237, B => n22044, S => n23067, Z => n5049
                           );
   U16636 : MUX2_X1 port map( A => n24239, B => n22046, S => n23067, Z => n5048
                           );
   U16637 : MUX2_X1 port map( A => n24241, B => n22048, S => n23067, Z => n5047
                           );
   U16638 : MUX2_X1 port map( A => n24243, B => n22050, S => n23068, Z => n5046
                           );
   U16639 : MUX2_X1 port map( A => n24245, B => n22161, S => n23068, Z => n5045
                           );
   U16640 : MUX2_X1 port map( A => n24247, B => n22163, S => n23068, Z => n5044
                           );
   U16641 : MUX2_X1 port map( A => n24249, B => n22052, S => n23068, Z => n5043
                           );
   U16642 : MUX2_X1 port map( A => n24251, B => n22166, S => n23068, Z => n5042
                           );
   U16643 : MUX2_X1 port map( A => n24253, B => n22167, S => n23068, Z => n5041
                           );
   U16644 : MUX2_X1 port map( A => n24255, B => n22169, S => n23068, Z => n5040
                           );
   U16645 : MUX2_X1 port map( A => n24257, B => n22171, S => n23068, Z => n5039
                           );
   U16646 : MUX2_X1 port map( A => n24259, B => n22054, S => n23068, Z => n5038
                           );
   U16647 : MUX2_X1 port map( A => n24261, B => n22174, S => n23068, Z => n5037
                           );
   U16648 : MUX2_X1 port map( A => n24263, B => n22176, S => n23068, Z => n5036
                           );
   U16649 : MUX2_X1 port map( A => n24265, B => n22177, S => n23068, Z => n5035
                           );
   U16650 : MUX2_X1 port map( A => n24267, B => n22178, S => n23069, Z => n5034
                           );
   U16651 : MUX2_X1 port map( A => n24269, B => n22180, S => n23069, Z => n5033
                           );
   U16652 : MUX2_X1 port map( A => n24271, B => n22181, S => n23069, Z => n5032
                           );
   U16653 : MUX2_X1 port map( A => n24273, B => n22183, S => n23069, Z => n5031
                           );
   U16654 : NAND3_X1 port map( A1 => N78, A2 => n22694, A3 => n24179, ZN => 
                           n24177);
   U16655 : NAND3_X1 port map( A1 => n22547, A2 => n22695, A3 => n24138, ZN => 
                           n24186);
   U16656 : OAI221_X1 port map( B1 => n24297, B2 => n24177, C1 => n24295, C2 =>
                           n24186, A => n23284, ZN => n24139);
   U16657 : INV_X1 port map( A => n24139, ZN => n24140);
   U16658 : MUX2_X1 port map( A => n24286, B => n22336, S => n23072, Z => n4582
                           );
   U16659 : MUX2_X1 port map( A => n24272, B => n22397, S => n23072, Z => n4581
                           );
   U16660 : MUX2_X1 port map( A => n24270, B => n22337, S => n23072, Z => n4580
                           );
   U16661 : MUX2_X1 port map( A => n24268, B => n22358, S => n23072, Z => n4579
                           );
   U16662 : MUX2_X1 port map( A => n24266, B => n22338, S => n23072, Z => n4578
                           );
   U16663 : MUX2_X1 port map( A => n24264, B => n22292, S => n23072, Z => n4577
                           );
   U16664 : MUX2_X1 port map( A => n24262, B => n22293, S => n23072, Z => n4576
                           );
   U16665 : MUX2_X1 port map( A => n24260, B => n22294, S => n23072, Z => n4575
                           );
   U16666 : MUX2_X1 port map( A => n24258, B => n22295, S => n23072, Z => n4574
                           );
   U16667 : MUX2_X1 port map( A => n24256, B => n22296, S => n23072, Z => n4573
                           );
   U16668 : MUX2_X1 port map( A => n24254, B => n22339, S => n23072, Z => n4572
                           );
   U16669 : MUX2_X1 port map( A => n24252, B => n22340, S => n23072, Z => n4571
                           );
   U16670 : MUX2_X1 port map( A => n24250, B => n22341, S => n23073, Z => n4570
                           );
   U16671 : MUX2_X1 port map( A => n24248, B => n22342, S => n23073, Z => n4569
                           );
   U16672 : MUX2_X1 port map( A => n24246, B => n22380, S => n23073, Z => n4568
                           );
   U16673 : MUX2_X1 port map( A => n24244, B => n22359, S => n23073, Z => n4567
                           );
   U16674 : MUX2_X1 port map( A => n24242, B => n22343, S => n23073, Z => n4566
                           );
   U16675 : MUX2_X1 port map( A => n24240, B => n22297, S => n23073, Z => n4565
                           );
   U16676 : MUX2_X1 port map( A => n24238, B => n22298, S => n23073, Z => n4564
                           );
   U16677 : MUX2_X1 port map( A => n24236, B => n22299, S => n23073, Z => n4563
                           );
   U16678 : MUX2_X1 port map( A => n24234, B => n22300, S => n23073, Z => n4562
                           );
   U16679 : MUX2_X1 port map( A => n24232, B => n22344, S => n23073, Z => n4561
                           );
   U16680 : MUX2_X1 port map( A => n24230, B => n22398, S => n23073, Z => n4560
                           );
   U16681 : MUX2_X1 port map( A => n24228, B => n22399, S => n23073, Z => n4559
                           );
   U16682 : MUX2_X1 port map( A => n24226, B => n22348, S => n23074, Z => n4558
                           );
   U16683 : MUX2_X1 port map( A => n24224, B => n22349, S => n23074, Z => n4557
                           );
   U16684 : MUX2_X1 port map( A => n24222, B => n22350, S => n23074, Z => n4556
                           );
   U16685 : MUX2_X1 port map( A => n24220, B => n22351, S => n23074, Z => n4555
                           );
   U16686 : MUX2_X1 port map( A => n24218, B => n22301, S => n23074, Z => n4554
                           );
   U16687 : MUX2_X1 port map( A => n24216, B => n22352, S => n23074, Z => n4553
                           );
   U16688 : MUX2_X1 port map( A => n24214, B => n22345, S => n23074, Z => n4552
                           );
   U16689 : MUX2_X1 port map( A => n24212, B => n22302, S => n23074, Z => n4551
                           );
   U16690 : MUX2_X1 port map( A => n24211, B => n22290, S => n23074, Z => n4550
                           );
   U16691 : MUX2_X1 port map( A => n24213, B => n22303, S => n23074, Z => n4549
                           );
   U16692 : MUX2_X1 port map( A => n24215, B => n22304, S => n23074, Z => n4548
                           );
   U16693 : MUX2_X1 port map( A => n24217, B => n22353, S => n23074, Z => n4547
                           );
   U16694 : MUX2_X1 port map( A => n24219, B => n22354, S => n23075, Z => n4546
                           );
   U16695 : MUX2_X1 port map( A => n24221, B => n22360, S => n23075, Z => n4545
                           );
   U16696 : MUX2_X1 port map( A => n24223, B => n22355, S => n23075, Z => n4544
                           );
   U16697 : MUX2_X1 port map( A => n24225, B => n22356, S => n23075, Z => n4543
                           );
   U16698 : MUX2_X1 port map( A => n24227, B => n22357, S => n23075, Z => n4542
                           );
   U16699 : MUX2_X1 port map( A => n24229, B => n22305, S => n23075, Z => n4541
                           );
   U16700 : MUX2_X1 port map( A => n24231, B => n22306, S => n23075, Z => n4540
                           );
   U16701 : MUX2_X1 port map( A => n24233, B => n22482, S => n23075, Z => n4539
                           );
   U16702 : MUX2_X1 port map( A => n24235, B => n22346, S => n23075, Z => n4538
                           );
   U16703 : MUX2_X1 port map( A => n24237, B => n22361, S => n23075, Z => n4537
                           );
   U16704 : MUX2_X1 port map( A => n24239, B => n22362, S => n23075, Z => n4536
                           );
   U16705 : MUX2_X1 port map( A => n24241, B => n22400, S => n23075, Z => n4535
                           );
   U16706 : MUX2_X1 port map( A => n24243, B => n22363, S => n23076, Z => n4534
                           );
   U16707 : MUX2_X1 port map( A => n24245, B => n22364, S => n23076, Z => n4533
                           );
   U16708 : MUX2_X1 port map( A => n24247, B => n22381, S => n23076, Z => n4532
                           );
   U16709 : MUX2_X1 port map( A => n24249, B => n22365, S => n23076, Z => n4531
                           );
   U16710 : MUX2_X1 port map( A => n24251, B => n22347, S => n23076, Z => n4530
                           );
   U16711 : MUX2_X1 port map( A => n24253, B => n22307, S => n23076, Z => n4529
                           );
   U16712 : MUX2_X1 port map( A => n24255, B => n22308, S => n23076, Z => n4528
                           );
   U16713 : MUX2_X1 port map( A => n24257, B => n22309, S => n23076, Z => n4527
                           );
   U16714 : MUX2_X1 port map( A => n24259, B => n22310, S => n23076, Z => n4526
                           );
   U16715 : MUX2_X1 port map( A => n24261, B => n22366, S => n23076, Z => n4525
                           );
   U16716 : MUX2_X1 port map( A => n24263, B => n22368, S => n23076, Z => n4524
                           );
   U16717 : MUX2_X1 port map( A => n24265, B => n22369, S => n23076, Z => n4523
                           );
   U16718 : MUX2_X1 port map( A => n24267, B => n22401, S => n23077, Z => n4522
                           );
   U16719 : MUX2_X1 port map( A => n24269, B => n22370, S => n23077, Z => n4521
                           );
   U16720 : MUX2_X1 port map( A => n24271, B => n22410, S => n23077, Z => n4520
                           );
   U16721 : MUX2_X1 port map( A => n24273, B => n22371, S => n23077, Z => n4519
                           );
   U16722 : NAND2_X1 port map( A1 => n22490, A2 => N76, ZN => n24294);
   U16723 : NAND2_X1 port map( A1 => n22532, A2 => n22688, ZN => n24291);
   U16724 : OAI221_X1 port map( B1 => n24294, B2 => n24177, C1 => n24291, C2 =>
                           n24186, A => n23284, ZN => n24141);
   U16725 : INV_X1 port map( A => n24141, ZN => n24142);
   U16726 : MUX2_X1 port map( A => n24286, B => n22373, S => n23080, Z => n4454
                           );
   U16727 : MUX2_X1 port map( A => n24272, B => n22374, S => n23080, Z => n4453
                           );
   U16728 : MUX2_X1 port map( A => n24270, B => n22375, S => n23080, Z => n4452
                           );
   U16729 : MUX2_X1 port map( A => n24268, B => n22376, S => n23080, Z => n4451
                           );
   U16730 : MUX2_X1 port map( A => n24266, B => n22367, S => n23080, Z => n4450
                           );
   U16731 : MUX2_X1 port map( A => n24264, B => n22311, S => n23080, Z => n4449
                           );
   U16732 : MUX2_X1 port map( A => n24262, B => n22312, S => n23080, Z => n4448
                           );
   U16733 : MUX2_X1 port map( A => n24260, B => n22313, S => n23080, Z => n4447
                           );
   U16734 : MUX2_X1 port map( A => n24258, B => n22314, S => n23080, Z => n4446
                           );
   U16735 : MUX2_X1 port map( A => n24256, B => n22315, S => n23080, Z => n4445
                           );
   U16736 : MUX2_X1 port map( A => n24254, B => n22377, S => n23080, Z => n4444
                           );
   U16737 : MUX2_X1 port map( A => n24252, B => n22382, S => n23080, Z => n4443
                           );
   U16738 : MUX2_X1 port map( A => n24250, B => n22383, S => n23081, Z => n4442
                           );
   U16739 : MUX2_X1 port map( A => n24248, B => n22384, S => n23081, Z => n4441
                           );
   U16740 : MUX2_X1 port map( A => n24246, B => n22385, S => n23081, Z => n4440
                           );
   U16741 : MUX2_X1 port map( A => n24244, B => n22386, S => n23081, Z => n4439
                           );
   U16742 : MUX2_X1 port map( A => n24242, B => n22316, S => n23081, Z => n4438
                           );
   U16743 : MUX2_X1 port map( A => n24240, B => n22317, S => n23081, Z => n4437
                           );
   U16744 : MUX2_X1 port map( A => n24238, B => n22318, S => n23081, Z => n4436
                           );
   U16745 : MUX2_X1 port map( A => n24236, B => n22319, S => n23081, Z => n4435
                           );
   U16746 : MUX2_X1 port map( A => n24234, B => n22320, S => n23081, Z => n4434
                           );
   U16747 : MUX2_X1 port map( A => n24232, B => n22378, S => n23081, Z => n4433
                           );
   U16748 : MUX2_X1 port map( A => n24230, B => n22321, S => n23081, Z => n4432
                           );
   U16749 : MUX2_X1 port map( A => n24228, B => n22387, S => n23081, Z => n4431
                           );
   U16750 : MUX2_X1 port map( A => n24226, B => n22388, S => n23082, Z => n4430
                           );
   U16751 : MUX2_X1 port map( A => n24224, B => n22402, S => n23082, Z => n4429
                           );
   U16752 : MUX2_X1 port map( A => n24222, B => n22389, S => n23082, Z => n4428
                           );
   U16753 : MUX2_X1 port map( A => n24220, B => n22390, S => n23082, Z => n4427
                           );
   U16754 : MUX2_X1 port map( A => n24218, B => n22322, S => n23082, Z => n4426
                           );
   U16755 : MUX2_X1 port map( A => n24216, B => n22323, S => n23082, Z => n4425
                           );
   U16756 : MUX2_X1 port map( A => n24214, B => n22324, S => n23082, Z => n4424
                           );
   U16757 : MUX2_X1 port map( A => n24212, B => n22325, S => n23082, Z => n4423
                           );
   U16758 : MUX2_X1 port map( A => n24211, B => n22372, S => n23082, Z => n4422
                           );
   U16759 : MUX2_X1 port map( A => n24213, B => n22326, S => n23082, Z => n4421
                           );
   U16760 : MUX2_X1 port map( A => n24215, B => n22379, S => n23082, Z => n4420
                           );
   U16761 : MUX2_X1 port map( A => n24217, B => n22391, S => n23082, Z => n4419
                           );
   U16762 : MUX2_X1 port map( A => n24219, B => n22392, S => n23083, Z => n4418
                           );
   U16763 : MUX2_X1 port map( A => n24221, B => n22393, S => n23083, Z => n4417
                           );
   U16764 : MUX2_X1 port map( A => n24223, B => n22394, S => n23083, Z => n4416
                           );
   U16765 : MUX2_X1 port map( A => n24225, B => n22395, S => n23083, Z => n4415
                           );
   U16766 : MUX2_X1 port map( A => n24227, B => n22327, S => n23083, Z => n4414
                           );
   U16767 : MUX2_X1 port map( A => n24229, B => n22328, S => n23083, Z => n4413
                           );
   U16768 : MUX2_X1 port map( A => n24231, B => n22329, S => n23083, Z => n4412
                           );
   U16769 : MUX2_X1 port map( A => n24233, B => n22483, S => n23083, Z => n4411
                           );
   U16770 : MUX2_X1 port map( A => n24235, B => n22330, S => n23083, Z => n4410
                           );
   U16771 : MUX2_X1 port map( A => n24237, B => n22396, S => n23083, Z => n4409
                           );
   U16772 : MUX2_X1 port map( A => n24239, B => n22403, S => n23083, Z => n4408
                           );
   U16773 : MUX2_X1 port map( A => n24241, B => n22404, S => n23083, Z => n4407
                           );
   U16774 : MUX2_X1 port map( A => n24243, B => n22405, S => n23084, Z => n4406
                           );
   U16775 : MUX2_X1 port map( A => n24245, B => n22406, S => n23084, Z => n4405
                           );
   U16776 : MUX2_X1 port map( A => n24247, B => n22407, S => n23084, Z => n4404
                           );
   U16777 : MUX2_X1 port map( A => n24249, B => n22408, S => n23084, Z => n4403
                           );
   U16778 : MUX2_X1 port map( A => n24251, B => n22331, S => n23084, Z => n4402
                           );
   U16779 : MUX2_X1 port map( A => n24253, B => n22332, S => n23084, Z => n4401
                           );
   U16780 : MUX2_X1 port map( A => n24255, B => n22333, S => n23084, Z => n4400
                           );
   U16781 : MUX2_X1 port map( A => n24257, B => n22334, S => n23084, Z => n4399
                           );
   U16782 : MUX2_X1 port map( A => n24259, B => n22335, S => n23084, Z => n4398
                           );
   U16783 : MUX2_X1 port map( A => n24261, B => n22409, S => n23084, Z => n4397
                           );
   U16784 : MUX2_X1 port map( A => n24263, B => n22411, S => n23084, Z => n4396
                           );
   U16785 : MUX2_X1 port map( A => n24265, B => n22412, S => n23084, Z => n4395
                           );
   U16786 : MUX2_X1 port map( A => n24267, B => n22413, S => n23085, Z => n4394
                           );
   U16787 : MUX2_X1 port map( A => n24269, B => n22414, S => n23085, Z => n4393
                           );
   U16788 : MUX2_X1 port map( A => n24271, B => n22415, S => n23085, Z => n4392
                           );
   U16789 : MUX2_X1 port map( A => n24273, B => n22416, S => n23085, Z => n4391
                           );
   U16790 : MUX2_X1 port map( A => n24143, B => CWP_2_port, S => n22768, Z => 
                           n24156);
   U16791 : NAND2_X1 port map( A1 => n22768, A2 => n24369, ZN => n24154);
   U16792 : INV_X1 port map( A => n24154, ZN => n24144);
   U16793 : MUX2_X1 port map( A => i_1_port, B => CWP_1_port, S => n22768, Z =>
                           n24151);
   U16794 : INV_X1 port map( A => n24151, ZN => n24146);
   U16795 : MUX2_X1 port map( A => i_0_port, B => CWP_0_port, S => n22768, Z =>
                           n24147);
   U16796 : OAI21_X1 port map( B1 => ADD_RD1(0), B2 => n20834, A => n24147, ZN 
                           => n24149);
   U16797 : INV_X1 port map( A => n24149, ZN => n24152);
   U16798 : OAI21_X1 port map( B1 => n24151, B2 => n24152, A => n22765, ZN => 
                           n24145);
   U16799 : OAI21_X1 port map( B1 => n24146, B2 => n24149, A => n24145, ZN => 
                           n24155);
   U16800 : INV_X1 port map( A => n24155, ZN => n24159);
   U16801 : INV_X1 port map( A => n24147, ZN => n24148);
   U16802 : NAND3_X1 port map( A1 => n22768, A2 => n24148, A3 => n24368, ZN => 
                           n24150);
   U16803 : NAND2_X1 port map( A1 => n24150, A2 => n24149, ZN => n18525);
   U16804 : XOR2_X1 port map( A => n24151, B => n22765, Z => n24153);
   U16805 : XOR2_X1 port map( A => n24153, B => n24152, Z => n25400);
   U16806 : INV_X1 port map( A => n25400, ZN => n18526);
   U16807 : INV_X1 port map( A => n18525, ZN => n25401);
   U16808 : INV_X1 port map( A => n24156, ZN => n24158);
   U16809 : OAI21_X1 port map( B1 => n24156, B2 => n24155, A => n24154, ZN => 
                           n24157);
   U16810 : OAI21_X1 port map( B1 => n24159, B2 => n24158, A => n24157, ZN => 
                           n24162);
   U16811 : INV_X1 port map( A => n24162, ZN => n24160);
   U16812 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => n22768, ZN => n24161);
   U16813 : NAND2_X1 port map( A1 => n24160, A2 => n24161, ZN => n24166);
   U16814 : INV_X1 port map( A => n24161, ZN => n24163);
   U16815 : NAND2_X1 port map( A1 => n24163, A2 => n24162, ZN => n24167);
   U16816 : NAND2_X1 port map( A1 => n24166, A2 => n24167, ZN => n24165);
   U16817 : MUX2_X1 port map( A => i_3_port, B => CWP_3_port, S => n22768, Z =>
                           n24164);
   U16818 : INV_X1 port map( A => n24164, ZN => n24168);
   U16819 : XOR2_X1 port map( A => n24165, B => n24168, Z => n24361);
   U16820 : INV_X1 port map( A => n24361, ZN => n24359);
   U16821 : INV_X1 port map( A => n24166, ZN => n24169);
   U16822 : OAI21_X1 port map( B1 => n24169, B2 => n24168, A => n24167, ZN => 
                           n24170);
   U16823 : XOR2_X1 port map( A => n24170, B => n3252, Z => n24172);
   U16824 : XOR2_X1 port map( A => n24170, B => n994, Z => n24171);
   U16825 : MUX2_X1 port map( A => n24172, B => n24171, S => n22768, Z => 
                           n24360);
   U16826 : INV_X1 port map( A => n24360, ZN => n24173);
   U16827 : NAND2_X1 port map( A1 => N76, A2 => n24176, ZN => n24300);
   U16828 : NAND2_X1 port map( A1 => n22688, A2 => n22796, ZN => n24298);
   U16829 : OAI221_X1 port map( B1 => n24300, B2 => n24177, C1 => n24298, C2 =>
                           n24186, A => n23284, ZN => n24174);
   U16830 : INV_X1 port map( A => n24174, ZN => n24274);
   U16831 : MUX2_X1 port map( A => n24211, B => n21284, S => n23088, Z => n4678
                           );
   U16832 : NAND2_X1 port map( A1 => n24176, A2 => n24175, ZN => n24305);
   U16833 : NAND3_X1 port map( A1 => n22506, A2 => n22497, A3 => n22797, ZN => 
                           n24302);
   U16834 : OAI221_X1 port map( B1 => n24305, B2 => n24177, C1 => n24302, C2 =>
                           n24186, A => n23284, ZN => n24178);
   U16835 : INV_X1 port map( A => n24178, ZN => n24275);
   U16836 : MUX2_X1 port map( A => n24211, B => n21841, S => n23096, Z => n4806
                           );
   U16837 : NAND3_X1 port map( A1 => N78, A2 => n22689, A3 => n24179, ZN => 
                           n24187);
   U16838 : OAI221_X1 port map( B1 => n24297, B2 => n24187, C1 => n24296, C2 =>
                           n24186, A => n23284, ZN => n24180);
   U16839 : INV_X1 port map( A => n24180, ZN => n24276);
   U16840 : MUX2_X1 port map( A => n24211, B => n22225, S => n23104, Z => n4614
                           );
   U16841 : NAND3_X1 port map( A1 => n22532, A2 => n22498, A3 => n22505, ZN => 
                           n24293);
   U16842 : OAI221_X1 port map( B1 => n24294, B2 => n24187, C1 => n24293, C2 =>
                           n24186, A => n23284, ZN => n24181);
   U16843 : INV_X1 port map( A => n24181, ZN => n24277);
   U16844 : MUX2_X1 port map( A => n24211, B => n22417, S => n23112, Z => n4486
                           );
   U16845 : NAND3_X1 port map( A1 => n22498, A2 => n22505, A3 => n22797, ZN => 
                           n24299);
   U16846 : OAI221_X1 port map( B1 => n24300, B2 => n24187, C1 => n24299, C2 =>
                           n24186, A => n23284, ZN => n24182);
   U16847 : INV_X1 port map( A => n24182, ZN => n24278);
   U16848 : MUX2_X1 port map( A => n24211, B => n21286, S => n23120, Z => n4742
                           );
   U16849 : NAND3_X1 port map( A1 => n22505, A2 => n22497, A3 => n22796, ZN => 
                           n24303);
   U16850 : OAI221_X1 port map( B1 => n24305, B2 => n24187, C1 => n24303, C2 =>
                           n24186, A => n23284, ZN => n24188);
   U16851 : INV_X1 port map( A => n24188, ZN => n24279);
   U16852 : MUX2_X1 port map( A => n24211, B => n21840, S => n23128, Z => n4870
                           );
   U16853 : OAI221_X1 port map( B1 => n24291, B2 => n24198, C1 => n24294, C2 =>
                           n24190, A => n23284, ZN => n24189);
   U16854 : INV_X1 port map( A => n24189, ZN => n24280);
   U16855 : MUX2_X1 port map( A => n24211, B => n21766, S => n23136, Z => n4934
                           );
   U16856 : INV_X1 port map( A => n24190, ZN => n24194);
   U16857 : INV_X1 port map( A => n24300, ZN => n24191);
   U16858 : AOI21_X1 port map( B1 => n24194, B2 => n24191, A => n16683, ZN => 
                           n24192);
   U16859 : OAI211_X1 port map( C1 => n24298, C2 => n24198, A => n23285, B => 
                           n24192, ZN => n24193);
   U16860 : INV_X1 port map( A => n24193, ZN => n24281);
   U16861 : MUX2_X1 port map( A => n24211, B => n20962, S => n23144, Z => n5190
                           );
   U16862 : INV_X1 port map( A => n24305, ZN => n24206);
   U16863 : AOI21_X1 port map( B1 => n24194, B2 => n24206, A => n16673, ZN => 
                           n24195);
   U16864 : OAI211_X1 port map( C1 => n24302, C2 => n24198, A => n23285, B => 
                           n24195, ZN => n24196);
   U16865 : INV_X1 port map( A => n24196, ZN => n24282);
   U16866 : MUX2_X1 port map( A => n24211, B => n21843, S => n23152, Z => n5318
                           );
   U16867 : OAI221_X1 port map( B1 => n24294, B2 => n24203, C1 => n24293, C2 =>
                           n24198, A => n23284, ZN => n24197);
   U16868 : INV_X1 port map( A => n24197, ZN => n24283);
   U16869 : MUX2_X1 port map( A => n24211, B => n22452, S => n23160, Z => n4998
                           );
   U16870 : INV_X1 port map( A => n24198, ZN => n24205);
   U16871 : INV_X1 port map( A => n24299, ZN => n24199);
   U16872 : AOI21_X1 port map( B1 => n24205, B2 => n24199, A => n16678, ZN => 
                           n24200);
   U16873 : OAI211_X1 port map( C1 => n24300, C2 => n24203, A => n23284, B => 
                           n24200, ZN => n24201);
   U16874 : INV_X1 port map( A => n24201, ZN => n24284);
   U16875 : MUX2_X1 port map( A => n24211, B => n21285, S => n23168, Z => n5254
                           );
   U16876 : NAND3_X1 port map( A1 => n24307, A2 => n24202, A3 => n22485, ZN => 
                           n16668);
   U16877 : INV_X1 port map( A => n24203, ZN => n24207);
   U16878 : INV_X1 port map( A => n24303, ZN => n24204);
   U16879 : AOI22_X1 port map( A1 => n24207, A2 => n24206, B1 => n24205, B2 => 
                           n24204, ZN => n24208);
   U16880 : OAI211_X1 port map( C1 => n16668, C2 => n24209, A => n23285, B => 
                           n24208, ZN => n24210);
   U16881 : INV_X1 port map( A => n24210, ZN => n24285);
   U16882 : MUX2_X1 port map( A => n24211, B => n21842, S => n23176, Z => n5382
                           );
   U16883 : MUX2_X1 port map( A => n24212, B => n21094, S => n23088, Z => n4679
                           );
   U16884 : MUX2_X1 port map( A => n24212, B => n21523, S => n23096, Z => n4807
                           );
   U16885 : MUX2_X1 port map( A => n24212, B => n22058, S => n23104, Z => n4615
                           );
   U16886 : MUX2_X1 port map( A => n24212, B => n22087, S => n23112, Z => n4487
                           );
   U16887 : MUX2_X1 port map( A => n24212, B => n21151, S => n23120, Z => n4743
                           );
   U16888 : MUX2_X1 port map( A => n24212, B => n21579, S => n23128, Z => n4871
                           );
   U16889 : MUX2_X1 port map( A => n24212, B => n21826, S => n23136, Z => n4935
                           );
   U16890 : MUX2_X1 port map( A => n24212, B => n20900, S => n23144, Z => n5191
                           );
   U16891 : MUX2_X1 port map( A => n24212, B => n21640, S => n23152, Z => n5319
                           );
   U16892 : MUX2_X1 port map( A => n24212, B => n22418, S => n23160, Z => n4999
                           );
   U16893 : MUX2_X1 port map( A => n24212, B => n21210, S => n23168, Z => n5255
                           );
   U16894 : MUX2_X1 port map( A => n24212, B => n21695, S => n23176, Z => n5383
                           );
   U16895 : MUX2_X1 port map( A => n24213, B => n21109, S => n23088, Z => n4677
                           );
   U16896 : MUX2_X1 port map( A => n24213, B => n21538, S => n23096, Z => n4805
                           );
   U16897 : MUX2_X1 port map( A => n24213, B => n22190, S => n23104, Z => n4613
                           );
   U16898 : MUX2_X1 port map( A => n24213, B => n22088, S => n23112, Z => n4485
                           );
   U16899 : MUX2_X1 port map( A => n24213, B => n21182, S => n23120, Z => n4741
                           );
   U16900 : MUX2_X1 port map( A => n24213, B => n21594, S => n23128, Z => n4869
                           );
   U16901 : MUX2_X1 port map( A => n24213, B => n21827, S => n23136, Z => n4933
                           );
   U16902 : MUX2_X1 port map( A => n24213, B => n20914, S => n23144, Z => n5189
                           );
   U16903 : MUX2_X1 port map( A => n24213, B => n21654, S => n23152, Z => n5317
                           );
   U16904 : MUX2_X1 port map( A => n24213, B => n22419, S => n23160, Z => n4997
                           );
   U16905 : MUX2_X1 port map( A => n24213, B => n21225, S => n23168, Z => n5253
                           );
   U16906 : MUX2_X1 port map( A => n24213, B => n21710, S => n23176, Z => n5381
                           );
   U16907 : MUX2_X1 port map( A => n24214, B => n21110, S => n23088, Z => n4680
                           );
   U16908 : MUX2_X1 port map( A => n24214, B => n21539, S => n23096, Z => n4808
                           );
   U16909 : MUX2_X1 port map( A => n24214, B => n22059, S => n23104, Z => n4616
                           );
   U16910 : MUX2_X1 port map( A => n24214, B => n22089, S => n23112, Z => n4488
                           );
   U16911 : MUX2_X1 port map( A => n24214, B => n21158, S => n23120, Z => n4744
                           );
   U16912 : MUX2_X1 port map( A => n24214, B => n21595, S => n23128, Z => n4872
                           );
   U16913 : MUX2_X1 port map( A => n24214, B => n21828, S => n23136, Z => n4936
                           );
   U16914 : MUX2_X1 port map( A => n24214, B => n20915, S => n23144, Z => n5192
                           );
   U16915 : MUX2_X1 port map( A => n24214, B => n21655, S => n23152, Z => n5320
                           );
   U16916 : MUX2_X1 port map( A => n24214, B => n22420, S => n23160, Z => n5000
                           );
   U16917 : MUX2_X1 port map( A => n24214, B => n21226, S => n23168, Z => n5256
                           );
   U16918 : MUX2_X1 port map( A => n24214, B => n21711, S => n23176, Z => n5384
                           );
   U16919 : MUX2_X1 port map( A => n24215, B => n21111, S => n23088, Z => n4676
                           );
   U16920 : MUX2_X1 port map( A => n24215, B => n21540, S => n23096, Z => n4804
                           );
   U16921 : MUX2_X1 port map( A => n24215, B => n22191, S => n23104, Z => n4612
                           );
   U16922 : MUX2_X1 port map( A => n24215, B => n22090, S => n23112, Z => n4484
                           );
   U16923 : MUX2_X1 port map( A => n24215, B => n21183, S => n23120, Z => n4740
                           );
   U16924 : MUX2_X1 port map( A => n24215, B => n21596, S => n23128, Z => n4868
                           );
   U16925 : MUX2_X1 port map( A => n24215, B => n21829, S => n23136, Z => n4932
                           );
   U16926 : MUX2_X1 port map( A => n24215, B => n20916, S => n23144, Z => n5188
                           );
   U16927 : MUX2_X1 port map( A => n24215, B => n21656, S => n23152, Z => n5316
                           );
   U16928 : MUX2_X1 port map( A => n24215, B => n22421, S => n23160, Z => n4996
                           );
   U16929 : MUX2_X1 port map( A => n24215, B => n21227, S => n23168, Z => n5252
                           );
   U16930 : MUX2_X1 port map( A => n24215, B => n21712, S => n23176, Z => n5380
                           );
   U16931 : MUX2_X1 port map( A => n24216, B => n21095, S => n23088, Z => n4681
                           );
   U16932 : MUX2_X1 port map( A => n24216, B => n21524, S => n23096, Z => n4809
                           );
   U16933 : MUX2_X1 port map( A => n24216, B => n22192, S => n23104, Z => n4617
                           );
   U16934 : MUX2_X1 port map( A => n24216, B => n22091, S => n23112, Z => n4489
                           );
   U16935 : MUX2_X1 port map( A => n24216, B => n21174, S => n23120, Z => n4745
                           );
   U16936 : MUX2_X1 port map( A => n24216, B => n21580, S => n23128, Z => n4873
                           );
   U16937 : MUX2_X1 port map( A => n24216, B => n21767, S => n23136, Z => n4937
                           );
   U16938 : MUX2_X1 port map( A => n24216, B => n20901, S => n23144, Z => n5193
                           );
   U16939 : MUX2_X1 port map( A => n24216, B => n21641, S => n23152, Z => n5321
                           );
   U16940 : MUX2_X1 port map( A => n24216, B => n22422, S => n23160, Z => n5001
                           );
   U16941 : MUX2_X1 port map( A => n24216, B => n21211, S => n23168, Z => n5257
                           );
   U16942 : MUX2_X1 port map( A => n24216, B => n21696, S => n23176, Z => n5385
                           );
   U16943 : MUX2_X1 port map( A => n24217, B => n21112, S => n23088, Z => n4675
                           );
   U16944 : MUX2_X1 port map( A => n24217, B => n21541, S => n23096, Z => n4803
                           );
   U16945 : MUX2_X1 port map( A => n24217, B => n22193, S => n23104, Z => n4611
                           );
   U16946 : MUX2_X1 port map( A => n24217, B => n22092, S => n23112, Z => n4483
                           );
   U16947 : MUX2_X1 port map( A => n24217, B => n21184, S => n23120, Z => n4739
                           );
   U16948 : MUX2_X1 port map( A => n24217, B => n21597, S => n23128, Z => n4867
                           );
   U16949 : MUX2_X1 port map( A => n24217, B => n21768, S => n23136, Z => n4931
                           );
   U16950 : MUX2_X1 port map( A => n24217, B => n20917, S => n23144, Z => n5187
                           );
   U16951 : MUX2_X1 port map( A => n24217, B => n21657, S => n23152, Z => n5315
                           );
   U16952 : MUX2_X1 port map( A => n24217, B => n22453, S => n23160, Z => n4995
                           );
   U16953 : MUX2_X1 port map( A => n24217, B => n21228, S => n23168, Z => n5251
                           );
   U16954 : MUX2_X1 port map( A => n24217, B => n21713, S => n23176, Z => n5379
                           );
   U16955 : MUX2_X1 port map( A => n24218, B => n21126, S => n23088, Z => n4682
                           );
   U16956 : MUX2_X1 port map( A => n24218, B => n21555, S => n23096, Z => n4810
                           );
   U16957 : MUX2_X1 port map( A => n24218, B => n22060, S => n23104, Z => n4618
                           );
   U16958 : MUX2_X1 port map( A => n24218, B => n22093, S => n23112, Z => n4490
                           );
   U16959 : MUX2_X1 port map( A => n24218, B => n21164, S => n23120, Z => n4746
                           );
   U16960 : MUX2_X1 port map( A => n24218, B => n21611, S => n23128, Z => n4874
                           );
   U16961 : MUX2_X1 port map( A => n24218, B => n21769, S => n23136, Z => n4938
                           );
   U16962 : MUX2_X1 port map( A => n24218, B => n20932, S => n23144, Z => n5194
                           );
   U16963 : MUX2_X1 port map( A => n24218, B => n21672, S => n23152, Z => n5322
                           );
   U16964 : MUX2_X1 port map( A => n24218, B => n22423, S => n23160, Z => n5002
                           );
   U16965 : MUX2_X1 port map( A => n24218, B => n21244, S => n23168, Z => n5258
                           );
   U16966 : MUX2_X1 port map( A => n24218, B => n21728, S => n23176, Z => n5386
                           );
   U16967 : MUX2_X1 port map( A => n24219, B => n21127, S => n23088, Z => n4674
                           );
   U16968 : MUX2_X1 port map( A => n24219, B => n21556, S => n23096, Z => n4802
                           );
   U16969 : MUX2_X1 port map( A => n24219, B => n22194, S => n23104, Z => n4610
                           );
   U16970 : MUX2_X1 port map( A => n24219, B => n22094, S => n23112, Z => n4482
                           );
   U16971 : MUX2_X1 port map( A => n24219, B => n21193, S => n23120, Z => n4738
                           );
   U16972 : MUX2_X1 port map( A => n24219, B => n21612, S => n23128, Z => n4866
                           );
   U16973 : MUX2_X1 port map( A => n24219, B => n21770, S => n23136, Z => n4930
                           );
   U16974 : MUX2_X1 port map( A => n24219, B => n20933, S => n23144, Z => n5186
                           );
   U16975 : MUX2_X1 port map( A => n24219, B => n21673, S => n23152, Z => n5314
                           );
   U16976 : MUX2_X1 port map( A => n24219, B => n22454, S => n23160, Z => n4994
                           );
   U16977 : MUX2_X1 port map( A => n24219, B => n21245, S => n23168, Z => n5250
                           );
   U16978 : MUX2_X1 port map( A => n24219, B => n21729, S => n23176, Z => n5378
                           );
   U16979 : MUX2_X1 port map( A => n24220, B => n21150, S => n23088, Z => n4683
                           );
   U16980 : MUX2_X1 port map( A => n24220, B => n21631, S => n23096, Z => n4811
                           );
   U16981 : MUX2_X1 port map( A => n24220, B => n22195, S => n23104, Z => n4619
                           );
   U16982 : MUX2_X1 port map( A => n24220, B => n22184, S => n23112, Z => n4491
                           );
   U16983 : MUX2_X1 port map( A => n24220, B => n21207, S => n23120, Z => n4747
                           );
   U16984 : MUX2_X1 port map( A => n24220, B => n21636, S => n23128, Z => n4875
                           );
   U16985 : MUX2_X1 port map( A => n24220, B => n21771, S => n23136, Z => n4939
                           );
   U16986 : MUX2_X1 port map( A => n24220, B => n20955, S => n23144, Z => n5195
                           );
   U16987 : MUX2_X1 port map( A => n24220, B => n21751, S => n23152, Z => n5323
                           );
   U16988 : MUX2_X1 port map( A => n24220, B => n22455, S => n23160, Z => n5003
                           );
   U16989 : MUX2_X1 port map( A => n24220, B => n21266, S => n23168, Z => n5259
                           );
   U16990 : MUX2_X1 port map( A => n24220, B => n21754, S => n23176, Z => n5387
                           );
   U16991 : MUX2_X1 port map( A => n24221, B => n21128, S => n23088, Z => n4673
                           );
   U16992 : MUX2_X1 port map( A => n24221, B => n21557, S => n23096, Z => n4801
                           );
   U16993 : MUX2_X1 port map( A => n24221, B => n22061, S => n23104, Z => n4609
                           );
   U16994 : MUX2_X1 port map( A => n24221, B => n22095, S => n23112, Z => n4481
                           );
   U16995 : MUX2_X1 port map( A => n24221, B => n21165, S => n23120, Z => n4737
                           );
   U16996 : MUX2_X1 port map( A => n24221, B => n21613, S => n23128, Z => n4865
                           );
   U16997 : MUX2_X1 port map( A => n24221, B => n21772, S => n23136, Z => n4929
                           );
   U16998 : MUX2_X1 port map( A => n24221, B => n20934, S => n23144, Z => n5185
                           );
   U16999 : MUX2_X1 port map( A => n24221, B => n21674, S => n23152, Z => n5313
                           );
   U17000 : MUX2_X1 port map( A => n24221, B => n22456, S => n23160, Z => n4993
                           );
   U17001 : MUX2_X1 port map( A => n24221, B => n21246, S => n23168, Z => n5249
                           );
   U17002 : MUX2_X1 port map( A => n24221, B => n21730, S => n23176, Z => n5377
                           );
   U17003 : MUX2_X1 port map( A => n24222, B => n21113, S => n23088, Z => n4684
                           );
   U17004 : MUX2_X1 port map( A => n24222, B => n21542, S => n23096, Z => n4812
                           );
   U17005 : MUX2_X1 port map( A => n24222, B => n22062, S => n23104, Z => n4620
                           );
   U17006 : MUX2_X1 port map( A => n24222, B => n22096, S => n23112, Z => n4492
                           );
   U17007 : MUX2_X1 port map( A => n24222, B => n21159, S => n23120, Z => n4748
                           );
   U17008 : MUX2_X1 port map( A => n24222, B => n21598, S => n23128, Z => n4876
                           );
   U17009 : MUX2_X1 port map( A => n24222, B => n21773, S => n23136, Z => n4940
                           );
   U17010 : MUX2_X1 port map( A => n24222, B => n20918, S => n23144, Z => n5196
                           );
   U17011 : MUX2_X1 port map( A => n24222, B => n21658, S => n23152, Z => n5324
                           );
   U17012 : MUX2_X1 port map( A => n24222, B => n22457, S => n23160, Z => n5004
                           );
   U17013 : MUX2_X1 port map( A => n24222, B => n21229, S => n23168, Z => n5260
                           );
   U17014 : MUX2_X1 port map( A => n24222, B => n21714, S => n23176, Z => n5388
                           );
   U17015 : MUX2_X1 port map( A => n24223, B => n21114, S => n23089, Z => n4672
                           );
   U17016 : MUX2_X1 port map( A => n24223, B => n21543, S => n23097, Z => n4800
                           );
   U17017 : MUX2_X1 port map( A => n24223, B => n22196, S => n23105, Z => n4608
                           );
   U17018 : MUX2_X1 port map( A => n24223, B => n22097, S => n23113, Z => n4480
                           );
   U17019 : MUX2_X1 port map( A => n24223, B => n21185, S => n23121, Z => n4736
                           );
   U17020 : MUX2_X1 port map( A => n24223, B => n21599, S => n23129, Z => n4864
                           );
   U17021 : MUX2_X1 port map( A => n24223, B => n21774, S => n23137, Z => n4928
                           );
   U17022 : MUX2_X1 port map( A => n24223, B => n20919, S => n23145, Z => n5184
                           );
   U17023 : MUX2_X1 port map( A => n24223, B => n21659, S => n23153, Z => n5312
                           );
   U17024 : MUX2_X1 port map( A => n24223, B => n22458, S => n23161, Z => n4992
                           );
   U17025 : MUX2_X1 port map( A => n24223, B => n21230, S => n23169, Z => n5248
                           );
   U17026 : MUX2_X1 port map( A => n24223, B => n21715, S => n23177, Z => n5376
                           );
   U17027 : MUX2_X1 port map( A => n24224, B => n21129, S => n23089, Z => n4685
                           );
   U17028 : MUX2_X1 port map( A => n24224, B => n21558, S => n23097, Z => n4813
                           );
   U17029 : MUX2_X1 port map( A => n24224, B => n22197, S => n23105, Z => n4621
                           );
   U17030 : MUX2_X1 port map( A => n24224, B => n22098, S => n23113, Z => n4493
                           );
   U17031 : MUX2_X1 port map( A => n24224, B => n21194, S => n23121, Z => n4749
                           );
   U17032 : MUX2_X1 port map( A => n24224, B => n21614, S => n23129, Z => n4877
                           );
   U17033 : MUX2_X1 port map( A => n24224, B => n21775, S => n23137, Z => n4941
                           );
   U17034 : MUX2_X1 port map( A => n24224, B => n20935, S => n23145, Z => n5197
                           );
   U17035 : MUX2_X1 port map( A => n24224, B => n21675, S => n23153, Z => n5325
                           );
   U17036 : MUX2_X1 port map( A => n24224, B => n22459, S => n23161, Z => n5005
                           );
   U17037 : MUX2_X1 port map( A => n24224, B => n21247, S => n23169, Z => n5261
                           );
   U17038 : MUX2_X1 port map( A => n24224, B => n21731, S => n23177, Z => n5389
                           );
   U17039 : MUX2_X1 port map( A => n24225, B => n21115, S => n23089, Z => n4671
                           );
   U17040 : MUX2_X1 port map( A => n24225, B => n21544, S => n23097, Z => n4799
                           );
   U17041 : MUX2_X1 port map( A => n24225, B => n22198, S => n23105, Z => n4607
                           );
   U17042 : MUX2_X1 port map( A => n24225, B => n22099, S => n23113, Z => n4479
                           );
   U17043 : MUX2_X1 port map( A => n24225, B => n21186, S => n23121, Z => n4735
                           );
   U17044 : MUX2_X1 port map( A => n24225, B => n21600, S => n23129, Z => n4863
                           );
   U17045 : MUX2_X1 port map( A => n24225, B => n21776, S => n23137, Z => n4927
                           );
   U17046 : MUX2_X1 port map( A => n24225, B => n20920, S => n23145, Z => n5183
                           );
   U17047 : MUX2_X1 port map( A => n24225, B => n21660, S => n23153, Z => n5311
                           );
   U17048 : MUX2_X1 port map( A => n24225, B => n22424, S => n23161, Z => n4991
                           );
   U17049 : MUX2_X1 port map( A => n24225, B => n21231, S => n23169, Z => n5247
                           );
   U17050 : MUX2_X1 port map( A => n24225, B => n21716, S => n23177, Z => n5375
                           );
   U17051 : MUX2_X1 port map( A => n24226, B => n21267, S => n23089, Z => n4686
                           );
   U17052 : MUX2_X1 port map( A => n24226, B => n21752, S => n23097, Z => n4814
                           );
   U17053 : MUX2_X1 port map( A => n24226, B => n22199, S => n23105, Z => n4622
                           );
   U17054 : MUX2_X1 port map( A => n24226, B => n22185, S => n23113, Z => n4494
                           );
   U17055 : MUX2_X1 port map( A => n24226, B => n21278, S => n23121, Z => n4750
                           );
   U17056 : MUX2_X1 port map( A => n24226, B => n21758, S => n23129, Z => n4878
                           );
   U17057 : MUX2_X1 port map( A => n24226, B => n21777, S => n23137, Z => n4942
                           );
   U17058 : MUX2_X1 port map( A => n24226, B => n20957, S => n23145, Z => n5198
                           );
   U17059 : MUX2_X1 port map( A => n24226, B => n21830, S => n23153, Z => n5326
                           );
   U17060 : MUX2_X1 port map( A => n24226, B => n22460, S => n23161, Z => n5006
                           );
   U17061 : MUX2_X1 port map( A => n24226, B => n21279, S => n23169, Z => n5262
                           );
   U17062 : MUX2_X1 port map( A => n24226, B => n21835, S => n23177, Z => n5390
                           );
   U17063 : MUX2_X1 port map( A => n24227, B => n21116, S => n23089, Z => n4670
                           );
   U17064 : MUX2_X1 port map( A => n24227, B => n21545, S => n23097, Z => n4798
                           );
   U17065 : MUX2_X1 port map( A => n24227, B => n22200, S => n23105, Z => n4606
                           );
   U17066 : MUX2_X1 port map( A => n24227, B => n22100, S => n23113, Z => n4478
                           );
   U17067 : MUX2_X1 port map( A => n24227, B => n21187, S => n23121, Z => n4734
                           );
   U17068 : MUX2_X1 port map( A => n24227, B => n21601, S => n23129, Z => n4862
                           );
   U17069 : MUX2_X1 port map( A => n24227, B => n21778, S => n23137, Z => n4926
                           );
   U17070 : MUX2_X1 port map( A => n24227, B => n20921, S => n23145, Z => n5182
                           );
   U17071 : MUX2_X1 port map( A => n24227, B => n21661, S => n23153, Z => n5310
                           );
   U17072 : MUX2_X1 port map( A => n24227, B => n22425, S => n23161, Z => n4990
                           );
   U17073 : MUX2_X1 port map( A => n24227, B => n21232, S => n23169, Z => n5246
                           );
   U17074 : MUX2_X1 port map( A => n24227, B => n21717, S => n23177, Z => n5374
                           );
   U17075 : MUX2_X1 port map( A => n24228, B => n21130, S => n23089, Z => n4687
                           );
   U17076 : MUX2_X1 port map( A => n24228, B => n21559, S => n23097, Z => n4815
                           );
   U17077 : MUX2_X1 port map( A => n24228, B => n22063, S => n23105, Z => n4623
                           );
   U17078 : MUX2_X1 port map( A => n24228, B => n22101, S => n23113, Z => n4495
                           );
   U17079 : MUX2_X1 port map( A => n24228, B => n21166, S => n23121, Z => n4751
                           );
   U17080 : MUX2_X1 port map( A => n24228, B => n21615, S => n23129, Z => n4879
                           );
   U17081 : MUX2_X1 port map( A => n24228, B => n21779, S => n23137, Z => n4943
                           );
   U17082 : MUX2_X1 port map( A => n24228, B => n20936, S => n23145, Z => n5199
                           );
   U17083 : MUX2_X1 port map( A => n24228, B => n21676, S => n23153, Z => n5327
                           );
   U17084 : MUX2_X1 port map( A => n24228, B => n22461, S => n23161, Z => n5007
                           );
   U17085 : MUX2_X1 port map( A => n24228, B => n21248, S => n23169, Z => n5263
                           );
   U17086 : MUX2_X1 port map( A => n24228, B => n21732, S => n23177, Z => n5391
                           );
   U17087 : MUX2_X1 port map( A => n24229, B => n21117, S => n23089, Z => n4669
                           );
   U17088 : MUX2_X1 port map( A => n24229, B => n21546, S => n23097, Z => n4797
                           );
   U17089 : MUX2_X1 port map( A => n24229, B => n22064, S => n23105, Z => n4605
                           );
   U17090 : MUX2_X1 port map( A => n24229, B => n22102, S => n23113, Z => n4477
                           );
   U17091 : MUX2_X1 port map( A => n24229, B => n21160, S => n23121, Z => n4733
                           );
   U17092 : MUX2_X1 port map( A => n24229, B => n21602, S => n23129, Z => n4861
                           );
   U17093 : MUX2_X1 port map( A => n24229, B => n21780, S => n23137, Z => n4925
                           );
   U17094 : MUX2_X1 port map( A => n24229, B => n20922, S => n23145, Z => n5181
                           );
   U17095 : MUX2_X1 port map( A => n24229, B => n21662, S => n23153, Z => n5309
                           );
   U17096 : MUX2_X1 port map( A => n24229, B => n22426, S => n23161, Z => n4989
                           );
   U17097 : MUX2_X1 port map( A => n24229, B => n21233, S => n23169, Z => n5245
                           );
   U17098 : MUX2_X1 port map( A => n24229, B => n21718, S => n23177, Z => n5373
                           );
   U17099 : MUX2_X1 port map( A => n24230, B => n21096, S => n23089, Z => n4688
                           );
   U17100 : MUX2_X1 port map( A => n24230, B => n21525, S => n23097, Z => n4816
                           );
   U17101 : MUX2_X1 port map( A => n24230, B => n22065, S => n23105, Z => n4624
                           );
   U17102 : MUX2_X1 port map( A => n24230, B => n22103, S => n23113, Z => n4496
                           );
   U17103 : MUX2_X1 port map( A => n24230, B => n21152, S => n23121, Z => n4752
                           );
   U17104 : MUX2_X1 port map( A => n24230, B => n21581, S => n23129, Z => n4880
                           );
   U17105 : MUX2_X1 port map( A => n24230, B => n21781, S => n23137, Z => n4944
                           );
   U17106 : MUX2_X1 port map( A => n24230, B => n20902, S => n23145, Z => n5200
                           );
   U17107 : MUX2_X1 port map( A => n24230, B => n21642, S => n23153, Z => n5328
                           );
   U17108 : MUX2_X1 port map( A => n24230, B => n22427, S => n23161, Z => n5008
                           );
   U17109 : MUX2_X1 port map( A => n24230, B => n21212, S => n23169, Z => n5264
                           );
   U17110 : MUX2_X1 port map( A => n24230, B => n21697, S => n23177, Z => n5392
                           );
   U17111 : MUX2_X1 port map( A => n24231, B => n21118, S => n23089, Z => n4668
                           );
   U17112 : MUX2_X1 port map( A => n24231, B => n21547, S => n23097, Z => n4796
                           );
   U17113 : MUX2_X1 port map( A => n24231, B => n22201, S => n23105, Z => n4604
                           );
   U17114 : MUX2_X1 port map( A => n24231, B => n22104, S => n23113, Z => n4476
                           );
   U17115 : MUX2_X1 port map( A => n24231, B => n21188, S => n23121, Z => n4732
                           );
   U17116 : MUX2_X1 port map( A => n24231, B => n21603, S => n23129, Z => n4860
                           );
   U17117 : MUX2_X1 port map( A => n24231, B => n21782, S => n23137, Z => n4924
                           );
   U17118 : MUX2_X1 port map( A => n24231, B => n20923, S => n23145, Z => n5180
                           );
   U17119 : MUX2_X1 port map( A => n24231, B => n21663, S => n23153, Z => n5308
                           );
   U17120 : MUX2_X1 port map( A => n24231, B => n22428, S => n23161, Z => n4988
                           );
   U17121 : MUX2_X1 port map( A => n24231, B => n21234, S => n23169, Z => n5244
                           );
   U17122 : MUX2_X1 port map( A => n24231, B => n21719, S => n23177, Z => n5372
                           );
   U17123 : MUX2_X1 port map( A => n24232, B => n21131, S => n23089, Z => n4689
                           );
   U17124 : MUX2_X1 port map( A => n24232, B => n21560, S => n23097, Z => n4817
                           );
   U17125 : MUX2_X1 port map( A => n24232, B => n22066, S => n23105, Z => n4625
                           );
   U17126 : MUX2_X1 port map( A => n24232, B => n22105, S => n23113, Z => n4497
                           );
   U17127 : MUX2_X1 port map( A => n24232, B => n21167, S => n23121, Z => n4753
                           );
   U17128 : MUX2_X1 port map( A => n24232, B => n21616, S => n23129, Z => n4881
                           );
   U17129 : MUX2_X1 port map( A => n24232, B => n21783, S => n23137, Z => n4945
                           );
   U17130 : MUX2_X1 port map( A => n24232, B => n20937, S => n23145, Z => n5201
                           );
   U17131 : MUX2_X1 port map( A => n24232, B => n21677, S => n23153, Z => n5329
                           );
   U17132 : MUX2_X1 port map( A => n24232, B => n22429, S => n23161, Z => n5009
                           );
   U17133 : MUX2_X1 port map( A => n24232, B => n21249, S => n23169, Z => n5265
                           );
   U17134 : MUX2_X1 port map( A => n24232, B => n21733, S => n23177, Z => n5393
                           );
   U17135 : MUX2_X1 port map( A => n24233, B => n21208, S => n23089, Z => n4667
                           );
   U17136 : MUX2_X1 port map( A => n24233, B => n21637, S => n23097, Z => n4795
                           );
   U17137 : MUX2_X1 port map( A => n24233, B => n22086, S => n23105, Z => n4603
                           );
   U17138 : MUX2_X1 port map( A => n24233, B => n22224, S => n23113, Z => n4475
                           );
   U17139 : MUX2_X1 port map( A => n24233, B => n21209, S => n23121, Z => n4731
                           );
   U17140 : MUX2_X1 port map( A => n24233, B => n21638, S => n23129, Z => n4859
                           );
   U17141 : MUX2_X1 port map( A => n24233, B => n21784, S => n23137, Z => n4923
                           );
   U17142 : MUX2_X1 port map( A => n24233, B => n20956, S => n23145, Z => n5179
                           );
   U17143 : MUX2_X1 port map( A => n24233, B => n21764, S => n23153, Z => n5307
                           );
   U17144 : MUX2_X1 port map( A => n24233, B => n22430, S => n23161, Z => n4987
                           );
   U17145 : MUX2_X1 port map( A => n24233, B => n21274, S => n23169, Z => n5243
                           );
   U17146 : MUX2_X1 port map( A => n24233, B => n21765, S => n23177, Z => n5371
                           );
   U17147 : MUX2_X1 port map( A => n24234, B => n21119, S => n23089, Z => n4690
                           );
   U17148 : MUX2_X1 port map( A => n24234, B => n21548, S => n23097, Z => n4818
                           );
   U17149 : MUX2_X1 port map( A => n24234, B => n22067, S => n23105, Z => n4626
                           );
   U17150 : MUX2_X1 port map( A => n24234, B => n22106, S => n23113, Z => n4498
                           );
   U17151 : MUX2_X1 port map( A => n24234, B => n21161, S => n23121, Z => n4754
                           );
   U17152 : MUX2_X1 port map( A => n24234, B => n21604, S => n23129, Z => n4882
                           );
   U17153 : MUX2_X1 port map( A => n24234, B => n21785, S => n23137, Z => n4946
                           );
   U17154 : MUX2_X1 port map( A => n24234, B => n20924, S => n23145, Z => n5202
                           );
   U17155 : MUX2_X1 port map( A => n24234, B => n21664, S => n23153, Z => n5330
                           );
   U17156 : MUX2_X1 port map( A => n24234, B => n22431, S => n23161, Z => n5010
                           );
   U17157 : MUX2_X1 port map( A => n24234, B => n21235, S => n23169, Z => n5266
                           );
   U17158 : MUX2_X1 port map( A => n24234, B => n21720, S => n23177, Z => n5394
                           );
   U17159 : MUX2_X1 port map( A => n24235, B => n21097, S => n23090, Z => n4666
                           );
   U17160 : MUX2_X1 port map( A => n24235, B => n21526, S => n23098, Z => n4794
                           );
   U17161 : MUX2_X1 port map( A => n24235, B => n22202, S => n23106, Z => n4602
                           );
   U17162 : MUX2_X1 port map( A => n24235, B => n22107, S => n23114, Z => n4474
                           );
   U17163 : MUX2_X1 port map( A => n24235, B => n21175, S => n23122, Z => n4730
                           );
   U17164 : MUX2_X1 port map( A => n24235, B => n21582, S => n23130, Z => n4858
                           );
   U17165 : MUX2_X1 port map( A => n24235, B => n21786, S => n23138, Z => n4922
                           );
   U17166 : MUX2_X1 port map( A => n24235, B => n20899, S => n23146, Z => n5178
                           );
   U17167 : MUX2_X1 port map( A => n24235, B => n21639, S => n23154, Z => n5306
                           );
   U17168 : MUX2_X1 port map( A => n24235, B => n22432, S => n23162, Z => n4986
                           );
   U17169 : MUX2_X1 port map( A => n24235, B => n21213, S => n23170, Z => n5242
                           );
   U17170 : MUX2_X1 port map( A => n24235, B => n21698, S => n23178, Z => n5370
                           );
   U17171 : MUX2_X1 port map( A => n24236, B => n21132, S => n23090, Z => n4691
                           );
   U17172 : MUX2_X1 port map( A => n24236, B => n21561, S => n23098, Z => n4819
                           );
   U17173 : MUX2_X1 port map( A => n24236, B => n22203, S => n23106, Z => n4627
                           );
   U17174 : MUX2_X1 port map( A => n24236, B => n22108, S => n23114, Z => n4499
                           );
   U17175 : MUX2_X1 port map( A => n24236, B => n21195, S => n23122, Z => n4755
                           );
   U17176 : MUX2_X1 port map( A => n24236, B => n21617, S => n23130, Z => n4883
                           );
   U17177 : MUX2_X1 port map( A => n24236, B => n21787, S => n23138, Z => n4947
                           );
   U17178 : MUX2_X1 port map( A => n24236, B => n20938, S => n23146, Z => n5203
                           );
   U17179 : MUX2_X1 port map( A => n24236, B => n21678, S => n23154, Z => n5331
                           );
   U17180 : MUX2_X1 port map( A => n24236, B => n22433, S => n23162, Z => n5011
                           );
   U17181 : MUX2_X1 port map( A => n24236, B => n21250, S => n23170, Z => n5267
                           );
   U17182 : MUX2_X1 port map( A => n24236, B => n21734, S => n23178, Z => n5395
                           );
   U17183 : MUX2_X1 port map( A => n24237, B => n21098, S => n23090, Z => n4665
                           );
   U17184 : MUX2_X1 port map( A => n24237, B => n21527, S => n23098, Z => n4793
                           );
   U17185 : MUX2_X1 port map( A => n24237, B => n22204, S => n23106, Z => n4601
                           );
   U17186 : MUX2_X1 port map( A => n24237, B => n22109, S => n23114, Z => n4473
                           );
   U17187 : MUX2_X1 port map( A => n24237, B => n21176, S => n23122, Z => n4729
                           );
   U17188 : MUX2_X1 port map( A => n24237, B => n21583, S => n23130, Z => n4857
                           );
   U17189 : MUX2_X1 port map( A => n24237, B => n21788, S => n23138, Z => n4921
                           );
   U17190 : MUX2_X1 port map( A => n24237, B => n20903, S => n23146, Z => n5177
                           );
   U17191 : MUX2_X1 port map( A => n24237, B => n21643, S => n23154, Z => n5305
                           );
   U17192 : MUX2_X1 port map( A => n24237, B => n22434, S => n23162, Z => n4985
                           );
   U17193 : MUX2_X1 port map( A => n24237, B => n21214, S => n23170, Z => n5241
                           );
   U17194 : MUX2_X1 port map( A => n24237, B => n21699, S => n23178, Z => n5369
                           );
   U17195 : MUX2_X1 port map( A => n24238, B => n21120, S => n23090, Z => n4692
                           );
   U17196 : MUX2_X1 port map( A => n24238, B => n21549, S => n23098, Z => n4820
                           );
   U17197 : MUX2_X1 port map( A => n24238, B => n22068, S => n23106, Z => n4628
                           );
   U17198 : MUX2_X1 port map( A => n24238, B => n22110, S => n23114, Z => n4500
                           );
   U17199 : MUX2_X1 port map( A => n24238, B => n21162, S => n23122, Z => n4756
                           );
   U17200 : MUX2_X1 port map( A => n24238, B => n21605, S => n23130, Z => n4884
                           );
   U17201 : MUX2_X1 port map( A => n24238, B => n21789, S => n23138, Z => n4948
                           );
   U17202 : MUX2_X1 port map( A => n24238, B => n20925, S => n23146, Z => n5204
                           );
   U17203 : MUX2_X1 port map( A => n24238, B => n21665, S => n23154, Z => n5332
                           );
   U17204 : MUX2_X1 port map( A => n24238, B => n22435, S => n23162, Z => n5012
                           );
   U17205 : MUX2_X1 port map( A => n24238, B => n21236, S => n23170, Z => n5268
                           );
   U17206 : MUX2_X1 port map( A => n24238, B => n21721, S => n23178, Z => n5396
                           );
   U17207 : MUX2_X1 port map( A => n24239, B => n21133, S => n23090, Z => n4664
                           );
   U17208 : MUX2_X1 port map( A => n24239, B => n21562, S => n23098, Z => n4792
                           );
   U17209 : MUX2_X1 port map( A => n24239, B => n22205, S => n23106, Z => n4600
                           );
   U17210 : MUX2_X1 port map( A => n24239, B => n22111, S => n23114, Z => n4472
                           );
   U17211 : MUX2_X1 port map( A => n24239, B => n21196, S => n23122, Z => n4728
                           );
   U17212 : MUX2_X1 port map( A => n24239, B => n21618, S => n23130, Z => n4856
                           );
   U17213 : MUX2_X1 port map( A => n24239, B => n21790, S => n23138, Z => n4920
                           );
   U17214 : MUX2_X1 port map( A => n24239, B => n20939, S => n23146, Z => n5176
                           );
   U17215 : MUX2_X1 port map( A => n24239, B => n21679, S => n23154, Z => n5304
                           );
   U17216 : MUX2_X1 port map( A => n24239, B => n22462, S => n23162, Z => n4984
                           );
   U17217 : MUX2_X1 port map( A => n24239, B => n21251, S => n23170, Z => n5240
                           );
   U17218 : MUX2_X1 port map( A => n24239, B => n21735, S => n23178, Z => n5368
                           );
   U17219 : MUX2_X1 port map( A => n24240, B => n21121, S => n23090, Z => n4693
                           );
   U17220 : MUX2_X1 port map( A => n24240, B => n21550, S => n23098, Z => n4821
                           );
   U17221 : MUX2_X1 port map( A => n24240, B => n22206, S => n23106, Z => n4629
                           );
   U17222 : MUX2_X1 port map( A => n24240, B => n22112, S => n23114, Z => n4501
                           );
   U17223 : MUX2_X1 port map( A => n24240, B => n21189, S => n23122, Z => n4757
                           );
   U17224 : MUX2_X1 port map( A => n24240, B => n21606, S => n23130, Z => n4885
                           );
   U17225 : MUX2_X1 port map( A => n24240, B => n21791, S => n23138, Z => n4949
                           );
   U17226 : MUX2_X1 port map( A => n24240, B => n20926, S => n23146, Z => n5205
                           );
   U17227 : MUX2_X1 port map( A => n24240, B => n21666, S => n23154, Z => n5333
                           );
   U17228 : MUX2_X1 port map( A => n24240, B => n22436, S => n23162, Z => n5013
                           );
   U17229 : MUX2_X1 port map( A => n24240, B => n21237, S => n23170, Z => n5269
                           );
   U17230 : MUX2_X1 port map( A => n24240, B => n21722, S => n23178, Z => n5397
                           );
   U17231 : MUX2_X1 port map( A => n24241, B => n21122, S => n23090, Z => n4663
                           );
   U17232 : MUX2_X1 port map( A => n24241, B => n21551, S => n23098, Z => n4791
                           );
   U17233 : MUX2_X1 port map( A => n24241, B => n22207, S => n23106, Z => n4599
                           );
   U17234 : MUX2_X1 port map( A => n24241, B => n22113, S => n23114, Z => n4471
                           );
   U17235 : MUX2_X1 port map( A => n24241, B => n21190, S => n23122, Z => n4727
                           );
   U17236 : MUX2_X1 port map( A => n24241, B => n21607, S => n23130, Z => n4855
                           );
   U17237 : MUX2_X1 port map( A => n24241, B => n21792, S => n23138, Z => n4919
                           );
   U17238 : MUX2_X1 port map( A => n24241, B => n20927, S => n23146, Z => n5175
                           );
   U17239 : MUX2_X1 port map( A => n24241, B => n21667, S => n23154, Z => n5303
                           );
   U17240 : MUX2_X1 port map( A => n24241, B => n22463, S => n23162, Z => n4983
                           );
   U17241 : MUX2_X1 port map( A => n24241, B => n21238, S => n23170, Z => n5239
                           );
   U17242 : MUX2_X1 port map( A => n24241, B => n21723, S => n23178, Z => n5367
                           );
   U17243 : MUX2_X1 port map( A => n24242, B => n21123, S => n23090, Z => n4694
                           );
   U17244 : MUX2_X1 port map( A => n24242, B => n21552, S => n23098, Z => n4822
                           );
   U17245 : MUX2_X1 port map( A => n24242, B => n22069, S => n23106, Z => n4630
                           );
   U17246 : MUX2_X1 port map( A => n24242, B => n22114, S => n23114, Z => n4502
                           );
   U17247 : MUX2_X1 port map( A => n24242, B => n21163, S => n23122, Z => n4758
                           );
   U17248 : MUX2_X1 port map( A => n24242, B => n21608, S => n23130, Z => n4886
                           );
   U17249 : MUX2_X1 port map( A => n24242, B => n21793, S => n23138, Z => n4950
                           );
   U17250 : MUX2_X1 port map( A => n24242, B => n20928, S => n23146, Z => n5206
                           );
   U17251 : MUX2_X1 port map( A => n24242, B => n21668, S => n23154, Z => n5334
                           );
   U17252 : MUX2_X1 port map( A => n24242, B => n22437, S => n23162, Z => n5014
                           );
   U17253 : MUX2_X1 port map( A => n24242, B => n21239, S => n23170, Z => n5270
                           );
   U17254 : MUX2_X1 port map( A => n24242, B => n21724, S => n23178, Z => n5398
                           );
   U17255 : MUX2_X1 port map( A => n24243, B => n21269, S => n23090, Z => n4662
                           );
   U17256 : MUX2_X1 port map( A => n24243, B => n21755, S => n23098, Z => n4790
                           );
   U17257 : MUX2_X1 port map( A => n24243, B => n22070, S => n23106, Z => n4598
                           );
   U17258 : MUX2_X1 port map( A => n24243, B => n22186, S => n23114, Z => n4470
                           );
   U17259 : MUX2_X1 port map( A => n24243, B => n21275, S => n23122, Z => n4726
                           );
   U17260 : MUX2_X1 port map( A => n24243, B => n21760, S => n23130, Z => n4854
                           );
   U17261 : MUX2_X1 port map( A => n24243, B => n21794, S => n23138, Z => n4918
                           );
   U17262 : MUX2_X1 port map( A => n24243, B => n20959, S => n23146, Z => n5174
                           );
   U17263 : MUX2_X1 port map( A => n24243, B => n21832, S => n23154, Z => n5302
                           );
   U17264 : MUX2_X1 port map( A => n24243, B => n22464, S => n23162, Z => n4982
                           );
   U17265 : MUX2_X1 port map( A => n24243, B => n21281, S => n23170, Z => n5238
                           );
   U17266 : MUX2_X1 port map( A => n24243, B => n21837, S => n23178, Z => n5366
                           );
   U17267 : MUX2_X1 port map( A => n24244, B => n21099, S => n23090, Z => n4695
                           );
   U17268 : MUX2_X1 port map( A => n24244, B => n21528, S => n23098, Z => n4823
                           );
   U17269 : MUX2_X1 port map( A => n24244, B => n22071, S => n23106, Z => n4631
                           );
   U17270 : MUX2_X1 port map( A => n24244, B => n22115, S => n23114, Z => n4503
                           );
   U17271 : MUX2_X1 port map( A => n24244, B => n21153, S => n23122, Z => n4759
                           );
   U17272 : MUX2_X1 port map( A => n24244, B => n21584, S => n23130, Z => n4887
                           );
   U17273 : MUX2_X1 port map( A => n24244, B => n21795, S => n23138, Z => n4951
                           );
   U17274 : MUX2_X1 port map( A => n24244, B => n20904, S => n23146, Z => n5207
                           );
   U17275 : MUX2_X1 port map( A => n24244, B => n21644, S => n23154, Z => n5335
                           );
   U17276 : MUX2_X1 port map( A => n24244, B => n22465, S => n23162, Z => n5015
                           );
   U17277 : MUX2_X1 port map( A => n24244, B => n21215, S => n23170, Z => n5271
                           );
   U17278 : MUX2_X1 port map( A => n24244, B => n21700, S => n23178, Z => n5399
                           );
   U17279 : MUX2_X1 port map( A => n24245, B => n21134, S => n23090, Z => n4661
                           );
   U17280 : MUX2_X1 port map( A => n24245, B => n21563, S => n23098, Z => n4789
                           );
   U17281 : MUX2_X1 port map( A => n24245, B => n22072, S => n23106, Z => n4597
                           );
   U17282 : MUX2_X1 port map( A => n24245, B => n22116, S => n23114, Z => n4469
                           );
   U17283 : MUX2_X1 port map( A => n24245, B => n21168, S => n23122, Z => n4725
                           );
   U17284 : MUX2_X1 port map( A => n24245, B => n21619, S => n23130, Z => n4853
                           );
   U17285 : MUX2_X1 port map( A => n24245, B => n21796, S => n23138, Z => n4917
                           );
   U17286 : MUX2_X1 port map( A => n24245, B => n20940, S => n23146, Z => n5173
                           );
   U17287 : MUX2_X1 port map( A => n24245, B => n21680, S => n23154, Z => n5301
                           );
   U17288 : MUX2_X1 port map( A => n24245, B => n22466, S => n23162, Z => n4981
                           );
   U17289 : MUX2_X1 port map( A => n24245, B => n21252, S => n23170, Z => n5237
                           );
   U17290 : MUX2_X1 port map( A => n24245, B => n21736, S => n23178, Z => n5365
                           );
   U17291 : MUX2_X1 port map( A => n24246, B => n21100, S => n23090, Z => n4696
                           );
   U17292 : MUX2_X1 port map( A => n24246, B => n21529, S => n23098, Z => n4824
                           );
   U17293 : MUX2_X1 port map( A => n24246, B => n22073, S => n23106, Z => n4632
                           );
   U17294 : MUX2_X1 port map( A => n24246, B => n22117, S => n23114, Z => n4504
                           );
   U17295 : MUX2_X1 port map( A => n24246, B => n21154, S => n23122, Z => n4760
                           );
   U17296 : MUX2_X1 port map( A => n24246, B => n21585, S => n23130, Z => n4888
                           );
   U17297 : MUX2_X1 port map( A => n24246, B => n21797, S => n23138, Z => n4952
                           );
   U17298 : MUX2_X1 port map( A => n24246, B => n20905, S => n23146, Z => n5208
                           );
   U17299 : MUX2_X1 port map( A => n24246, B => n21645, S => n23154, Z => n5336
                           );
   U17300 : MUX2_X1 port map( A => n24246, B => n22467, S => n23162, Z => n5016
                           );
   U17301 : MUX2_X1 port map( A => n24246, B => n21216, S => n23170, Z => n5272
                           );
   U17302 : MUX2_X1 port map( A => n24246, B => n21701, S => n23178, Z => n5400
                           );
   U17303 : MUX2_X1 port map( A => n24247, B => n21270, S => n23091, Z => n4660
                           );
   U17304 : MUX2_X1 port map( A => n24247, B => n21756, S => n23099, Z => n4788
                           );
   U17305 : MUX2_X1 port map( A => n24247, B => n22074, S => n23107, Z => n4596
                           );
   U17306 : MUX2_X1 port map( A => n24247, B => n22187, S => n23115, Z => n4468
                           );
   U17307 : MUX2_X1 port map( A => n24247, B => n21276, S => n23123, Z => n4724
                           );
   U17308 : MUX2_X1 port map( A => n24247, B => n21761, S => n23131, Z => n4852
                           );
   U17309 : MUX2_X1 port map( A => n24247, B => n21798, S => n23139, Z => n4916
                           );
   U17310 : MUX2_X1 port map( A => n24247, B => n20960, S => n23147, Z => n5172
                           );
   U17311 : MUX2_X1 port map( A => n24247, B => n21833, S => n23155, Z => n5300
                           );
   U17312 : MUX2_X1 port map( A => n24247, B => n22468, S => n23163, Z => n4980
                           );
   U17313 : MUX2_X1 port map( A => n24247, B => n21282, S => n23171, Z => n5236
                           );
   U17314 : MUX2_X1 port map( A => n24247, B => n21838, S => n23179, Z => n5364
                           );
   U17315 : MUX2_X1 port map( A => n24248, B => n21271, S => n23091, Z => n4697
                           );
   U17316 : MUX2_X1 port map( A => n24248, B => n21757, S => n23099, Z => n4825
                           );
   U17317 : MUX2_X1 port map( A => n24248, B => n22075, S => n23107, Z => n4633
                           );
   U17318 : MUX2_X1 port map( A => n24248, B => n22188, S => n23115, Z => n4505
                           );
   U17319 : MUX2_X1 port map( A => n24248, B => n21277, S => n23123, Z => n4761
                           );
   U17320 : MUX2_X1 port map( A => n24248, B => n21762, S => n23131, Z => n4889
                           );
   U17321 : MUX2_X1 port map( A => n24248, B => n21799, S => n23139, Z => n4953
                           );
   U17322 : MUX2_X1 port map( A => n24248, B => n20961, S => n23147, Z => n5209
                           );
   U17323 : MUX2_X1 port map( A => n24248, B => n21834, S => n23155, Z => n5337
                           );
   U17324 : MUX2_X1 port map( A => n24248, B => n22469, S => n23163, Z => n5017
                           );
   U17325 : MUX2_X1 port map( A => n24248, B => n21283, S => n23171, Z => n5273
                           );
   U17326 : MUX2_X1 port map( A => n24248, B => n21839, S => n23179, Z => n5401
                           );
   U17327 : MUX2_X1 port map( A => n24249, B => n21124, S => n23091, Z => n4659
                           );
   U17328 : MUX2_X1 port map( A => n24249, B => n21553, S => n23099, Z => n4787
                           );
   U17329 : MUX2_X1 port map( A => n24249, B => n22208, S => n23107, Z => n4595
                           );
   U17330 : MUX2_X1 port map( A => n24249, B => n22118, S => n23115, Z => n4467
                           );
   U17331 : MUX2_X1 port map( A => n24249, B => n21191, S => n23123, Z => n4723
                           );
   U17332 : MUX2_X1 port map( A => n24249, B => n21609, S => n23131, Z => n4851
                           );
   U17333 : MUX2_X1 port map( A => n24249, B => n21800, S => n23139, Z => n4915
                           );
   U17334 : MUX2_X1 port map( A => n24249, B => n20929, S => n23147, Z => n5171
                           );
   U17335 : MUX2_X1 port map( A => n24249, B => n21669, S => n23155, Z => n5299
                           );
   U17336 : MUX2_X1 port map( A => n24249, B => n22438, S => n23163, Z => n4979
                           );
   U17337 : MUX2_X1 port map( A => n24249, B => n21240, S => n23171, Z => n5235
                           );
   U17338 : MUX2_X1 port map( A => n24249, B => n21725, S => n23179, Z => n5363
                           );
   U17339 : MUX2_X1 port map( A => n24250, B => n21101, S => n23091, Z => n4698
                           );
   U17340 : MUX2_X1 port map( A => n24250, B => n21530, S => n23099, Z => n4826
                           );
   U17341 : MUX2_X1 port map( A => n24250, B => n22076, S => n23107, Z => n4634
                           );
   U17342 : MUX2_X1 port map( A => n24250, B => n22119, S => n23115, Z => n4506
                           );
   U17343 : MUX2_X1 port map( A => n24250, B => n21155, S => n23123, Z => n4762
                           );
   U17344 : MUX2_X1 port map( A => n24250, B => n21586, S => n23131, Z => n4890
                           );
   U17345 : MUX2_X1 port map( A => n24250, B => n21801, S => n23139, Z => n4954
                           );
   U17346 : MUX2_X1 port map( A => n24250, B => n20906, S => n23147, Z => n5210
                           );
   U17347 : MUX2_X1 port map( A => n24250, B => n21646, S => n23155, Z => n5338
                           );
   U17348 : MUX2_X1 port map( A => n24250, B => n22470, S => n23163, Z => n5018
                           );
   U17349 : MUX2_X1 port map( A => n24250, B => n21217, S => n23171, Z => n5274
                           );
   U17350 : MUX2_X1 port map( A => n24250, B => n21702, S => n23179, Z => n5402
                           );
   U17351 : MUX2_X1 port map( A => n24251, B => n21268, S => n23091, Z => n4658
                           );
   U17352 : MUX2_X1 port map( A => n24251, B => n21753, S => n23099, Z => n4786
                           );
   U17353 : MUX2_X1 port map( A => n24251, B => n22077, S => n23107, Z => n4594
                           );
   U17354 : MUX2_X1 port map( A => n24251, B => n22189, S => n23115, Z => n4466
                           );
   U17355 : MUX2_X1 port map( A => n24251, B => n21273, S => n23123, Z => n4722
                           );
   U17356 : MUX2_X1 port map( A => n24251, B => n21759, S => n23131, Z => n4850
                           );
   U17357 : MUX2_X1 port map( A => n24251, B => n21802, S => n23139, Z => n4914
                           );
   U17358 : MUX2_X1 port map( A => n24251, B => n20958, S => n23147, Z => n5170
                           );
   U17359 : MUX2_X1 port map( A => n24251, B => n21831, S => n23155, Z => n5298
                           );
   U17360 : MUX2_X1 port map( A => n24251, B => n22439, S => n23163, Z => n4978
                           );
   U17361 : MUX2_X1 port map( A => n24251, B => n21280, S => n23171, Z => n5234
                           );
   U17362 : MUX2_X1 port map( A => n24251, B => n21836, S => n23179, Z => n5362
                           );
   U17363 : MUX2_X1 port map( A => n24252, B => n21135, S => n23091, Z => n4699
                           );
   U17364 : MUX2_X1 port map( A => n24252, B => n21564, S => n23099, Z => n4827
                           );
   U17365 : MUX2_X1 port map( A => n24252, B => n22078, S => n23107, Z => n4635
                           );
   U17366 : MUX2_X1 port map( A => n24252, B => n22120, S => n23115, Z => n4507
                           );
   U17367 : MUX2_X1 port map( A => n24252, B => n21169, S => n23123, Z => n4763
                           );
   U17368 : MUX2_X1 port map( A => n24252, B => n21620, S => n23131, Z => n4891
                           );
   U17369 : MUX2_X1 port map( A => n24252, B => n21803, S => n23139, Z => n4955
                           );
   U17370 : MUX2_X1 port map( A => n24252, B => n20941, S => n23147, Z => n5211
                           );
   U17371 : MUX2_X1 port map( A => n24252, B => n21681, S => n23155, Z => n5339
                           );
   U17372 : MUX2_X1 port map( A => n24252, B => n22471, S => n23163, Z => n5019
                           );
   U17373 : MUX2_X1 port map( A => n24252, B => n21253, S => n23171, Z => n5275
                           );
   U17374 : MUX2_X1 port map( A => n24252, B => n21737, S => n23179, Z => n5403
                           );
   U17375 : MUX2_X1 port map( A => n24253, B => n21102, S => n23091, Z => n4657
                           );
   U17376 : MUX2_X1 port map( A => n24253, B => n21531, S => n23099, Z => n4785
                           );
   U17377 : MUX2_X1 port map( A => n24253, B => n22079, S => n23107, Z => n4593
                           );
   U17378 : MUX2_X1 port map( A => n24253, B => n22121, S => n23115, Z => n4465
                           );
   U17379 : MUX2_X1 port map( A => n24253, B => n21156, S => n23123, Z => n4721
                           );
   U17380 : MUX2_X1 port map( A => n24253, B => n21587, S => n23131, Z => n4849
                           );
   U17381 : MUX2_X1 port map( A => n24253, B => n21804, S => n23139, Z => n4913
                           );
   U17382 : MUX2_X1 port map( A => n24253, B => n20907, S => n23147, Z => n5169
                           );
   U17383 : MUX2_X1 port map( A => n24253, B => n21647, S => n23155, Z => n5297
                           );
   U17384 : MUX2_X1 port map( A => n24253, B => n22440, S => n23163, Z => n4977
                           );
   U17385 : MUX2_X1 port map( A => n24253, B => n21218, S => n23171, Z => n5233
                           );
   U17386 : MUX2_X1 port map( A => n24253, B => n21703, S => n23179, Z => n5361
                           );
   U17387 : MUX2_X1 port map( A => n24254, B => n21136, S => n23091, Z => n4700
                           );
   U17388 : MUX2_X1 port map( A => n24254, B => n21565, S => n23099, Z => n4828
                           );
   U17389 : MUX2_X1 port map( A => n24254, B => n22080, S => n23107, Z => n4636
                           );
   U17390 : MUX2_X1 port map( A => n24254, B => n22122, S => n23115, Z => n4508
                           );
   U17391 : MUX2_X1 port map( A => n24254, B => n21170, S => n23123, Z => n4764
                           );
   U17392 : MUX2_X1 port map( A => n24254, B => n21621, S => n23131, Z => n4892
                           );
   U17393 : MUX2_X1 port map( A => n24254, B => n21805, S => n23139, Z => n4956
                           );
   U17394 : MUX2_X1 port map( A => n24254, B => n20942, S => n23147, Z => n5212
                           );
   U17395 : MUX2_X1 port map( A => n24254, B => n21682, S => n23155, Z => n5340
                           );
   U17396 : MUX2_X1 port map( A => n24254, B => n22441, S => n23163, Z => n5020
                           );
   U17397 : MUX2_X1 port map( A => n24254, B => n21254, S => n23171, Z => n5276
                           );
   U17398 : MUX2_X1 port map( A => n24254, B => n21738, S => n23179, Z => n5404
                           );
   U17399 : MUX2_X1 port map( A => n24255, B => n21103, S => n23091, Z => n4656
                           );
   U17400 : MUX2_X1 port map( A => n24255, B => n21532, S => n23099, Z => n4784
                           );
   U17401 : MUX2_X1 port map( A => n24255, B => n22081, S => n23107, Z => n4592
                           );
   U17402 : MUX2_X1 port map( A => n24255, B => n22123, S => n23115, Z => n4464
                           );
   U17403 : MUX2_X1 port map( A => n24255, B => n21157, S => n23123, Z => n4720
                           );
   U17404 : MUX2_X1 port map( A => n24255, B => n21588, S => n23131, Z => n4848
                           );
   U17405 : MUX2_X1 port map( A => n24255, B => n21806, S => n23139, Z => n4912
                           );
   U17406 : MUX2_X1 port map( A => n24255, B => n20908, S => n23147, Z => n5168
                           );
   U17407 : MUX2_X1 port map( A => n24255, B => n21648, S => n23155, Z => n5296
                           );
   U17408 : MUX2_X1 port map( A => n24255, B => n22442, S => n23163, Z => n4976
                           );
   U17409 : MUX2_X1 port map( A => n24255, B => n21219, S => n23171, Z => n5232
                           );
   U17410 : MUX2_X1 port map( A => n24255, B => n21704, S => n23179, Z => n5360
                           );
   U17411 : MUX2_X1 port map( A => n24256, B => n21137, S => n23091, Z => n4701
                           );
   U17412 : MUX2_X1 port map( A => n24256, B => n21566, S => n23099, Z => n4829
                           );
   U17413 : MUX2_X1 port map( A => n24256, B => n22209, S => n23107, Z => n4637
                           );
   U17414 : MUX2_X1 port map( A => n24256, B => n22124, S => n23115, Z => n4509
                           );
   U17415 : MUX2_X1 port map( A => n24256, B => n21197, S => n23123, Z => n4765
                           );
   U17416 : MUX2_X1 port map( A => n24256, B => n21622, S => n23131, Z => n4893
                           );
   U17417 : MUX2_X1 port map( A => n24256, B => n21807, S => n23139, Z => n4957
                           );
   U17418 : MUX2_X1 port map( A => n24256, B => n20943, S => n23147, Z => n5213
                           );
   U17419 : MUX2_X1 port map( A => n24256, B => n21683, S => n23155, Z => n5341
                           );
   U17420 : MUX2_X1 port map( A => n24256, B => n22443, S => n23163, Z => n5021
                           );
   U17421 : MUX2_X1 port map( A => n24256, B => n21255, S => n23171, Z => n5277
                           );
   U17422 : MUX2_X1 port map( A => n24256, B => n21739, S => n23179, Z => n5405
                           );
   U17423 : MUX2_X1 port map( A => n24257, B => n21138, S => n23091, Z => n4655
                           );
   U17424 : MUX2_X1 port map( A => n24257, B => n21567, S => n23099, Z => n4783
                           );
   U17425 : MUX2_X1 port map( A => n24257, B => n22082, S => n23107, Z => n4591
                           );
   U17426 : MUX2_X1 port map( A => n24257, B => n22125, S => n23115, Z => n4463
                           );
   U17427 : MUX2_X1 port map( A => n24257, B => n21171, S => n23123, Z => n4719
                           );
   U17428 : MUX2_X1 port map( A => n24257, B => n21623, S => n23131, Z => n4847
                           );
   U17429 : MUX2_X1 port map( A => n24257, B => n21808, S => n23139, Z => n4911
                           );
   U17430 : MUX2_X1 port map( A => n24257, B => n20944, S => n23147, Z => n5167
                           );
   U17431 : MUX2_X1 port map( A => n24257, B => n21684, S => n23155, Z => n5295
                           );
   U17432 : MUX2_X1 port map( A => n24257, B => n22444, S => n23163, Z => n4975
                           );
   U17433 : MUX2_X1 port map( A => n24257, B => n21256, S => n23171, Z => n5231
                           );
   U17434 : MUX2_X1 port map( A => n24257, B => n21740, S => n23179, Z => n5359
                           );
   U17435 : MUX2_X1 port map( A => n24258, B => n21104, S => n23091, Z => n4702
                           );
   U17436 : MUX2_X1 port map( A => n24258, B => n21533, S => n23099, Z => n4830
                           );
   U17437 : MUX2_X1 port map( A => n24258, B => n22210, S => n23107, Z => n4638
                           );
   U17438 : MUX2_X1 port map( A => n24258, B => n22126, S => n23115, Z => n4510
                           );
   U17439 : MUX2_X1 port map( A => n24258, B => n21177, S => n23123, Z => n4766
                           );
   U17440 : MUX2_X1 port map( A => n24258, B => n21589, S => n23131, Z => n4894
                           );
   U17441 : MUX2_X1 port map( A => n24258, B => n21809, S => n23139, Z => n4958
                           );
   U17442 : MUX2_X1 port map( A => n24258, B => n20909, S => n23147, Z => n5214
                           );
   U17443 : MUX2_X1 port map( A => n24258, B => n21649, S => n23155, Z => n5342
                           );
   U17444 : MUX2_X1 port map( A => n24258, B => n22445, S => n23163, Z => n5022
                           );
   U17445 : MUX2_X1 port map( A => n24258, B => n21220, S => n23171, Z => n5278
                           );
   U17446 : MUX2_X1 port map( A => n24258, B => n21705, S => n23179, Z => n5406
                           );
   U17447 : MUX2_X1 port map( A => n24259, B => n21139, S => n23092, Z => n4654
                           );
   U17448 : MUX2_X1 port map( A => n24259, B => n21568, S => n23100, Z => n4782
                           );
   U17449 : MUX2_X1 port map( A => n24259, B => n22083, S => n23108, Z => n4590
                           );
   U17450 : MUX2_X1 port map( A => n24259, B => n22127, S => n23116, Z => n4462
                           );
   U17451 : MUX2_X1 port map( A => n24259, B => n21172, S => n23124, Z => n4718
                           );
   U17452 : MUX2_X1 port map( A => n24259, B => n21624, S => n23132, Z => n4846
                           );
   U17453 : MUX2_X1 port map( A => n24259, B => n21810, S => n23140, Z => n4910
                           );
   U17454 : MUX2_X1 port map( A => n24259, B => n20945, S => n23148, Z => n5166
                           );
   U17455 : MUX2_X1 port map( A => n24259, B => n21685, S => n23156, Z => n5294
                           );
   U17456 : MUX2_X1 port map( A => n24259, B => n22446, S => n23164, Z => n4974
                           );
   U17457 : MUX2_X1 port map( A => n24259, B => n21257, S => n23172, Z => n5230
                           );
   U17458 : MUX2_X1 port map( A => n24259, B => n21741, S => n23180, Z => n5358
                           );
   U17459 : MUX2_X1 port map( A => n24260, B => n21125, S => n23092, Z => n4703
                           );
   U17460 : MUX2_X1 port map( A => n24260, B => n21554, S => n23100, Z => n4831
                           );
   U17461 : MUX2_X1 port map( A => n24260, B => n22211, S => n23108, Z => n4639
                           );
   U17462 : MUX2_X1 port map( A => n24260, B => n22128, S => n23116, Z => n4511
                           );
   U17463 : MUX2_X1 port map( A => n24260, B => n21192, S => n23124, Z => n4767
                           );
   U17464 : MUX2_X1 port map( A => n24260, B => n21610, S => n23132, Z => n4895
                           );
   U17465 : MUX2_X1 port map( A => n24260, B => n21811, S => n23140, Z => n4959
                           );
   U17466 : MUX2_X1 port map( A => n24260, B => n20930, S => n23148, Z => n5215
                           );
   U17467 : MUX2_X1 port map( A => n24260, B => n21670, S => n23156, Z => n5343
                           );
   U17468 : MUX2_X1 port map( A => n24260, B => n22447, S => n23164, Z => n5023
                           );
   U17469 : MUX2_X1 port map( A => n24260, B => n21241, S => n23172, Z => n5279
                           );
   U17470 : MUX2_X1 port map( A => n24260, B => n21726, S => n23180, Z => n5407
                           );
   U17471 : MUX2_X1 port map( A => n24261, B => n21105, S => n23092, Z => n4653
                           );
   U17472 : MUX2_X1 port map( A => n24261, B => n21534, S => n23100, Z => n4781
                           );
   U17473 : MUX2_X1 port map( A => n24261, B => n22212, S => n23108, Z => n4589
                           );
   U17474 : MUX2_X1 port map( A => n24261, B => n22129, S => n23116, Z => n4461
                           );
   U17475 : MUX2_X1 port map( A => n24261, B => n21178, S => n23124, Z => n4717
                           );
   U17476 : MUX2_X1 port map( A => n24261, B => n21590, S => n23132, Z => n4845
                           );
   U17477 : MUX2_X1 port map( A => n24261, B => n21812, S => n23140, Z => n4909
                           );
   U17478 : MUX2_X1 port map( A => n24261, B => n20910, S => n23148, Z => n5165
                           );
   U17479 : MUX2_X1 port map( A => n24261, B => n21650, S => n23156, Z => n5293
                           );
   U17480 : MUX2_X1 port map( A => n24261, B => n22448, S => n23164, Z => n4973
                           );
   U17481 : MUX2_X1 port map( A => n24261, B => n21221, S => n23172, Z => n5229
                           );
   U17482 : MUX2_X1 port map( A => n24261, B => n21706, S => n23180, Z => n5357
                           );
   U17483 : MUX2_X1 port map( A => n24262, B => n21140, S => n23092, Z => n4704
                           );
   U17484 : MUX2_X1 port map( A => n24262, B => n21569, S => n23100, Z => n4832
                           );
   U17485 : MUX2_X1 port map( A => n24262, B => n22213, S => n23108, Z => n4640
                           );
   U17486 : MUX2_X1 port map( A => n24262, B => n22130, S => n23116, Z => n4512
                           );
   U17487 : MUX2_X1 port map( A => n24262, B => n21198, S => n23124, Z => n4768
                           );
   U17488 : MUX2_X1 port map( A => n24262, B => n21625, S => n23132, Z => n4896
                           );
   U17489 : MUX2_X1 port map( A => n24262, B => n21813, S => n23140, Z => n4960
                           );
   U17490 : MUX2_X1 port map( A => n24262, B => n20946, S => n23148, Z => n5216
                           );
   U17491 : MUX2_X1 port map( A => n24262, B => n21686, S => n23156, Z => n5344
                           );
   U17492 : MUX2_X1 port map( A => n24262, B => n22449, S => n23164, Z => n5024
                           );
   U17493 : MUX2_X1 port map( A => n24262, B => n21258, S => n23172, Z => n5280
                           );
   U17494 : MUX2_X1 port map( A => n24262, B => n21742, S => n23180, Z => n5408
                           );
   U17495 : MUX2_X1 port map( A => n24263, B => n21141, S => n23092, Z => n4652
                           );
   U17496 : MUX2_X1 port map( A => n24263, B => n21570, S => n23100, Z => n4780
                           );
   U17497 : MUX2_X1 port map( A => n24263, B => n22214, S => n23108, Z => n4588
                           );
   U17498 : MUX2_X1 port map( A => n24263, B => n22131, S => n23116, Z => n4460
                           );
   U17499 : MUX2_X1 port map( A => n24263, B => n21199, S => n23124, Z => n4716
                           );
   U17500 : MUX2_X1 port map( A => n24263, B => n21626, S => n23132, Z => n4844
                           );
   U17501 : MUX2_X1 port map( A => n24263, B => n21814, S => n23140, Z => n4908
                           );
   U17502 : MUX2_X1 port map( A => n24263, B => n20947, S => n23148, Z => n5164
                           );
   U17503 : MUX2_X1 port map( A => n24263, B => n21687, S => n23156, Z => n5292
                           );
   U17504 : MUX2_X1 port map( A => n24263, B => n22472, S => n23164, Z => n4972
                           );
   U17505 : MUX2_X1 port map( A => n24263, B => n21259, S => n23172, Z => n5228
                           );
   U17506 : MUX2_X1 port map( A => n24263, B => n21743, S => n23180, Z => n5356
                           );
   U17507 : MUX2_X1 port map( A => n24264, B => n21106, S => n23092, Z => n4705
                           );
   U17508 : MUX2_X1 port map( A => n24264, B => n21535, S => n23100, Z => n4833
                           );
   U17509 : MUX2_X1 port map( A => n24264, B => n22215, S => n23108, Z => n4641
                           );
   U17510 : MUX2_X1 port map( A => n24264, B => n22132, S => n23116, Z => n4513
                           );
   U17511 : MUX2_X1 port map( A => n24264, B => n21179, S => n23124, Z => n4769
                           );
   U17512 : MUX2_X1 port map( A => n24264, B => n21591, S => n23132, Z => n4897
                           );
   U17513 : MUX2_X1 port map( A => n24264, B => n21815, S => n23140, Z => n4961
                           );
   U17514 : MUX2_X1 port map( A => n24264, B => n20911, S => n23148, Z => n5217
                           );
   U17515 : MUX2_X1 port map( A => n24264, B => n21651, S => n23156, Z => n5345
                           );
   U17516 : MUX2_X1 port map( A => n24264, B => n22450, S => n23164, Z => n5025
                           );
   U17517 : MUX2_X1 port map( A => n24264, B => n21222, S => n23172, Z => n5281
                           );
   U17518 : MUX2_X1 port map( A => n24264, B => n21707, S => n23180, Z => n5409
                           );
   U17519 : MUX2_X1 port map( A => n24265, B => n21142, S => n23092, Z => n4651
                           );
   U17520 : MUX2_X1 port map( A => n24265, B => n21571, S => n23100, Z => n4779
                           );
   U17521 : MUX2_X1 port map( A => n24265, B => n22216, S => n23108, Z => n4587
                           );
   U17522 : MUX2_X1 port map( A => n24265, B => n22133, S => n23116, Z => n4459
                           );
   U17523 : MUX2_X1 port map( A => n24265, B => n21200, S => n23124, Z => n4715
                           );
   U17524 : MUX2_X1 port map( A => n24265, B => n21627, S => n23132, Z => n4843
                           );
   U17525 : MUX2_X1 port map( A => n24265, B => n21816, S => n23140, Z => n4907
                           );
   U17526 : MUX2_X1 port map( A => n24265, B => n20948, S => n23148, Z => n5163
                           );
   U17527 : MUX2_X1 port map( A => n24265, B => n21688, S => n23156, Z => n5291
                           );
   U17528 : MUX2_X1 port map( A => n24265, B => n22473, S => n23164, Z => n4971
                           );
   U17529 : MUX2_X1 port map( A => n24265, B => n21260, S => n23172, Z => n5227
                           );
   U17530 : MUX2_X1 port map( A => n24265, B => n21744, S => n23180, Z => n5355
                           );
   U17531 : MUX2_X1 port map( A => n24266, B => n21143, S => n23092, Z => n4706
                           );
   U17532 : MUX2_X1 port map( A => n24266, B => n21572, S => n23100, Z => n4834
                           );
   U17533 : MUX2_X1 port map( A => n24266, B => n22217, S => n23108, Z => n4642
                           );
   U17534 : MUX2_X1 port map( A => n24266, B => n22134, S => n23116, Z => n4514
                           );
   U17535 : MUX2_X1 port map( A => n24266, B => n21201, S => n23124, Z => n4770
                           );
   U17536 : MUX2_X1 port map( A => n24266, B => n21628, S => n23132, Z => n4898
                           );
   U17537 : MUX2_X1 port map( A => n24266, B => n21817, S => n23140, Z => n4962
                           );
   U17538 : MUX2_X1 port map( A => n24266, B => n20949, S => n23148, Z => n5218
                           );
   U17539 : MUX2_X1 port map( A => n24266, B => n21689, S => n23156, Z => n5346
                           );
   U17540 : MUX2_X1 port map( A => n24266, B => n22451, S => n23164, Z => n5026
                           );
   U17541 : MUX2_X1 port map( A => n24266, B => n21243, S => n23172, Z => n5282
                           );
   U17542 : MUX2_X1 port map( A => n24266, B => n21745, S => n23180, Z => n5410
                           );
   U17543 : MUX2_X1 port map( A => n24267, B => n21107, S => n23092, Z => n4650
                           );
   U17544 : MUX2_X1 port map( A => n24267, B => n21536, S => n23100, Z => n4778
                           );
   U17545 : MUX2_X1 port map( A => n24267, B => n22218, S => n23108, Z => n4586
                           );
   U17546 : MUX2_X1 port map( A => n24267, B => n22135, S => n23116, Z => n4458
                           );
   U17547 : MUX2_X1 port map( A => n24267, B => n21180, S => n23124, Z => n4714
                           );
   U17548 : MUX2_X1 port map( A => n24267, B => n21592, S => n23132, Z => n4842
                           );
   U17549 : MUX2_X1 port map( A => n24267, B => n21818, S => n23140, Z => n4906
                           );
   U17550 : MUX2_X1 port map( A => n24267, B => n20912, S => n23148, Z => n5162
                           );
   U17551 : MUX2_X1 port map( A => n24267, B => n21652, S => n23156, Z => n5290
                           );
   U17552 : MUX2_X1 port map( A => n24267, B => n22474, S => n23164, Z => n4970
                           );
   U17553 : MUX2_X1 port map( A => n24267, B => n21223, S => n23172, Z => n5226
                           );
   U17554 : MUX2_X1 port map( A => n24267, B => n21708, S => n23180, Z => n5354
                           );
   U17555 : MUX2_X1 port map( A => n24268, B => n21144, S => n23092, Z => n4707
                           );
   U17556 : MUX2_X1 port map( A => n24268, B => n21573, S => n23100, Z => n4835
                           );
   U17557 : MUX2_X1 port map( A => n24268, B => n22084, S => n23108, Z => n4643
                           );
   U17558 : MUX2_X1 port map( A => n24268, B => n22136, S => n23116, Z => n4515
                           );
   U17559 : MUX2_X1 port map( A => n24268, B => n21173, S => n23124, Z => n4771
                           );
   U17560 : MUX2_X1 port map( A => n24268, B => n21629, S => n23132, Z => n4899
                           );
   U17561 : MUX2_X1 port map( A => n24268, B => n21819, S => n23140, Z => n4963
                           );
   U17562 : MUX2_X1 port map( A => n24268, B => n20950, S => n23148, Z => n5219
                           );
   U17563 : MUX2_X1 port map( A => n24268, B => n21690, S => n23156, Z => n5347
                           );
   U17564 : MUX2_X1 port map( A => n24268, B => n22475, S => n23164, Z => n5027
                           );
   U17565 : MUX2_X1 port map( A => n24268, B => n21261, S => n23172, Z => n5283
                           );
   U17566 : MUX2_X1 port map( A => n24268, B => n21746, S => n23180, Z => n5411
                           );
   U17567 : MUX2_X1 port map( A => n24269, B => n21145, S => n23092, Z => n4649
                           );
   U17568 : MUX2_X1 port map( A => n24269, B => n21574, S => n23100, Z => n4777
                           );
   U17569 : MUX2_X1 port map( A => n24269, B => n22219, S => n23108, Z => n4585
                           );
   U17570 : MUX2_X1 port map( A => n24269, B => n22137, S => n23116, Z => n4457
                           );
   U17571 : MUX2_X1 port map( A => n24269, B => n21202, S => n23124, Z => n4713
                           );
   U17572 : MUX2_X1 port map( A => n24269, B => n21630, S => n23132, Z => n4841
                           );
   U17573 : MUX2_X1 port map( A => n24269, B => n21820, S => n23140, Z => n4905
                           );
   U17574 : MUX2_X1 port map( A => n24269, B => n20951, S => n23148, Z => n5161
                           );
   U17575 : MUX2_X1 port map( A => n24269, B => n21691, S => n23156, Z => n5289
                           );
   U17576 : MUX2_X1 port map( A => n24269, B => n22476, S => n23164, Z => n4969
                           );
   U17577 : MUX2_X1 port map( A => n24269, B => n21262, S => n23172, Z => n5225
                           );
   U17578 : MUX2_X1 port map( A => n24269, B => n21747, S => n23180, Z => n5353
                           );
   U17579 : MUX2_X1 port map( A => n24270, B => n21108, S => n23092, Z => n4708
                           );
   U17580 : MUX2_X1 port map( A => n24270, B => n21537, S => n23100, Z => n4836
                           );
   U17581 : MUX2_X1 port map( A => n24270, B => n22220, S => n23108, Z => n4644
                           );
   U17582 : MUX2_X1 port map( A => n24270, B => n22138, S => n23116, Z => n4516
                           );
   U17583 : MUX2_X1 port map( A => n24270, B => n21181, S => n23124, Z => n4772
                           );
   U17584 : MUX2_X1 port map( A => n24270, B => n21593, S => n23132, Z => n4900
                           );
   U17585 : MUX2_X1 port map( A => n24270, B => n21821, S => n23140, Z => n4964
                           );
   U17586 : MUX2_X1 port map( A => n24270, B => n20913, S => n23148, Z => n5220
                           );
   U17587 : MUX2_X1 port map( A => n24270, B => n21653, S => n23156, Z => n5348
                           );
   U17588 : MUX2_X1 port map( A => n24270, B => n22477, S => n23164, Z => n5028
                           );
   U17589 : MUX2_X1 port map( A => n24270, B => n21224, S => n23172, Z => n5284
                           );
   U17590 : MUX2_X1 port map( A => n24270, B => n21709, S => n23180, Z => n5412
                           );
   U17591 : MUX2_X1 port map( A => n24271, B => n21147, S => n23093, Z => n4648
                           );
   U17592 : MUX2_X1 port map( A => n24271, B => n21576, S => n23101, Z => n4776
                           );
   U17593 : MUX2_X1 port map( A => n24271, B => n22221, S => n23109, Z => n4584
                           );
   U17594 : MUX2_X1 port map( A => n24271, B => n22139, S => n23117, Z => n4456
                           );
   U17595 : MUX2_X1 port map( A => n24271, B => n21204, S => n23125, Z => n4712
                           );
   U17596 : MUX2_X1 port map( A => n24271, B => n21633, S => n23133, Z => n4840
                           );
   U17597 : MUX2_X1 port map( A => n24271, B => n21822, S => n23141, Z => n4904
                           );
   U17598 : MUX2_X1 port map( A => n24271, B => n20952, S => n23149, Z => n5160
                           );
   U17599 : MUX2_X1 port map( A => n24271, B => n21692, S => n23157, Z => n5288
                           );
   U17600 : MUX2_X1 port map( A => n24271, B => n22478, S => n23165, Z => n4968
                           );
   U17601 : MUX2_X1 port map( A => n24271, B => n21263, S => n23173, Z => n5224
                           );
   U17602 : MUX2_X1 port map( A => n24271, B => n21748, S => n23181, Z => n5352
                           );
   U17603 : MUX2_X1 port map( A => n24272, B => n21148, S => n23093, Z => n4709
                           );
   U17604 : MUX2_X1 port map( A => n24272, B => n21577, S => n23101, Z => n4837
                           );
   U17605 : MUX2_X1 port map( A => n24272, B => n22222, S => n23109, Z => n4645
                           );
   U17606 : MUX2_X1 port map( A => n24272, B => n22140, S => n23117, Z => n4517
                           );
   U17607 : MUX2_X1 port map( A => n24272, B => n21205, S => n23125, Z => n4773
                           );
   U17608 : MUX2_X1 port map( A => n24272, B => n21634, S => n23133, Z => n4901
                           );
   U17609 : MUX2_X1 port map( A => n24272, B => n21823, S => n23141, Z => n4965
                           );
   U17610 : MUX2_X1 port map( A => n24272, B => n20953, S => n23149, Z => n5221
                           );
   U17611 : MUX2_X1 port map( A => n24272, B => n21693, S => n23157, Z => n5349
                           );
   U17612 : MUX2_X1 port map( A => n24272, B => n22479, S => n23165, Z => n5029
                           );
   U17613 : MUX2_X1 port map( A => n24272, B => n21264, S => n23173, Z => n5285
                           );
   U17614 : MUX2_X1 port map( A => n24272, B => n21749, S => n23181, Z => n5413
                           );
   U17615 : MUX2_X1 port map( A => n24273, B => n21146, S => n23093, Z => n4647
                           );
   U17616 : MUX2_X1 port map( A => n24273, B => n21575, S => n23101, Z => n4775
                           );
   U17617 : MUX2_X1 port map( A => n24273, B => n22085, S => n23109, Z => n4583
                           );
   U17618 : MUX2_X1 port map( A => n24273, B => n22141, S => n23117, Z => n4455
                           );
   U17619 : MUX2_X1 port map( A => n24273, B => n21203, S => n23125, Z => n4711
                           );
   U17620 : MUX2_X1 port map( A => n24273, B => n21632, S => n23133, Z => n4839
                           );
   U17621 : MUX2_X1 port map( A => n24273, B => n21824, S => n23141, Z => n4903
                           );
   U17622 : MUX2_X1 port map( A => n24273, B => n20931, S => n23149, Z => n5159
                           );
   U17623 : MUX2_X1 port map( A => n24273, B => n21671, S => n23157, Z => n5287
                           );
   U17624 : MUX2_X1 port map( A => n24273, B => n22480, S => n23165, Z => n4967
                           );
   U17625 : MUX2_X1 port map( A => n24273, B => n21242, S => n23173, Z => n5223
                           );
   U17626 : MUX2_X1 port map( A => n24273, B => n21727, S => n23181, Z => n5351
                           );
   U17627 : MUX2_X1 port map( A => n24286, B => n21149, S => n23093, Z => n4710
                           );
   U17628 : MUX2_X1 port map( A => n24286, B => n21578, S => n23101, Z => n4838
                           );
   U17629 : MUX2_X1 port map( A => n24286, B => n22223, S => n23109, Z => n4646
                           );
   U17630 : MUX2_X1 port map( A => n24286, B => n22142, S => n23117, Z => n4518
                           );
   U17631 : MUX2_X1 port map( A => n24286, B => n21206, S => n23125, Z => n4774
                           );
   U17632 : MUX2_X1 port map( A => n24286, B => n21635, S => n23133, Z => n4902
                           );
   U17633 : MUX2_X1 port map( A => n24286, B => n21825, S => n23141, Z => n4966
                           );
   U17634 : MUX2_X1 port map( A => n24286, B => n20954, S => n23149, Z => n5222
                           );
   U17635 : MUX2_X1 port map( A => n24286, B => n21694, S => n23157, Z => n5350
                           );
   U17636 : MUX2_X1 port map( A => n24286, B => n22481, S => n23165, Z => n5030
                           );
   U17637 : MUX2_X1 port map( A => n24286, B => n21265, S => n23173, Z => n5286
                           );
   U17638 : MUX2_X1 port map( A => n24286, B => n21750, S => n23181, Z => n5414
                           );
   U17639 : NAND3_X1 port map( A1 => n22547, A2 => n22495, A3 => n22695, ZN => 
                           n24289);
   U17640 : NAND2_X1 port map( A1 => n22678, A2 => n22694, ZN => n24287);
   U17641 : OAI221_X1 port map( B1 => n24291, B2 => n24289, C1 => n24294, C2 =>
                           n24287, A => n23284, ZN => n16735);
   U17642 : NAND2_X1 port map( A1 => n22678, A2 => n22689, ZN => n24288);
   U17643 : OAI221_X1 port map( B1 => n24293, B2 => n24289, C1 => n24294, C2 =>
                           n24288, A => n23284, ZN => n16734);
   U17644 : OAI221_X1 port map( B1 => n24295, B2 => n24289, C1 => n24297, C2 =>
                           n24287, A => n23284, ZN => n16733);
   U17645 : OAI221_X1 port map( B1 => n24296, B2 => n24289, C1 => n24297, C2 =>
                           n24288, A => n23284, ZN => n16732);
   U17646 : OAI221_X1 port map( B1 => n24298, B2 => n24289, C1 => n24300, C2 =>
                           n24287, A => n23283, ZN => n16731);
   U17647 : OAI221_X1 port map( B1 => n24299, B2 => n24289, C1 => n24300, C2 =>
                           n24288, A => n23283, ZN => n16730);
   U17648 : OAI221_X1 port map( B1 => n24302, B2 => n24289, C1 => n24305, C2 =>
                           n24287, A => n23283, ZN => n16728);
   U17649 : OAI221_X1 port map( B1 => n24303, B2 => n24289, C1 => n24305, C2 =>
                           n24288, A => n23283, ZN => n16725);
   U17650 : NAND3_X1 port map( A1 => n22495, A2 => n22695, A3 => n24290, ZN => 
                           n24304);
   U17651 : NAND3_X1 port map( A1 => n22694, A2 => n22508, A3 => n24292, ZN => 
                           n24301);
   U17652 : OAI221_X1 port map( B1 => n24304, B2 => n24291, C1 => n24301, C2 =>
                           n24294, A => n23283, ZN => n16724);
   U17653 : NAND3_X1 port map( A1 => n22508, A2 => n22689, A3 => n24292, ZN => 
                           n24306);
   U17654 : OAI221_X1 port map( B1 => n24306, B2 => n24294, C1 => n24304, C2 =>
                           n24293, A => n23284, ZN => n16722);
   U17655 : OAI221_X1 port map( B1 => n24304, B2 => n24295, C1 => n24301, C2 =>
                           n24297, A => n23283, ZN => n16721);
   U17656 : OAI221_X1 port map( B1 => n24306, B2 => n24297, C1 => n24304, C2 =>
                           n24296, A => n23283, ZN => n16720);
   U17657 : OAI221_X1 port map( B1 => n24304, B2 => n24298, C1 => n24301, C2 =>
                           n24300, A => n23283, ZN => n16719);
   U17658 : OAI221_X1 port map( B1 => n24306, B2 => n24300, C1 => n24304, C2 =>
                           n24299, A => n23283, ZN => n16718);
   U17659 : OAI221_X1 port map( B1 => n24304, B2 => n24302, C1 => n24305, C2 =>
                           n24301, A => n23283, ZN => n16716);
   U17660 : OAI221_X1 port map( B1 => n24306, B2 => n24305, C1 => n24304, C2 =>
                           n24303, A => n23283, ZN => n16713);
   U17661 : NAND2_X1 port map( A1 => RD2, A2 => n24307, ZN => n16581);
   U17662 : MUX2_X1 port map( A => n18526, B => n25408, S => n22768, Z => 
                           n24324);
   U17663 : MUX2_X1 port map( A => n18525, B => n25409, S => n22768, Z => 
                           n24327);
   U17664 : OAI21_X1 port map( B1 => n3046, B2 => n24327, A => n3044, ZN => 
                           n24322);
   U17665 : INV_X1 port map( A => n24322, ZN => n24309);
   U17666 : INV_X1 port map( A => n24327, ZN => n24308);
   U17667 : NAND3_X1 port map( A1 => n24308, A2 => CWP_1_port, A3 => CWP_0_port
                           , ZN => n24323);
   U17668 : OAI21_X1 port map( B1 => n24324, B2 => n24309, A => n24323, ZN => 
                           n24313);
   U17669 : INV_X1 port map( A => n24313, ZN => n24329);
   U17670 : INV_X1 port map( A => n25402, ZN => n24311);
   U17671 : INV_X1 port map( A => ADD_RD2(2), ZN => n24310);
   U17672 : MUX2_X1 port map( A => n24311, B => n24310, S => n22768, Z => 
                           n24328);
   U17673 : OAI21_X1 port map( B1 => n3045, B2 => n24329, A => n24328, ZN => 
                           n24312);
   U17674 : OAI21_X1 port map( B1 => n24313, B2 => CWP_2_port, A => n24312, ZN 
                           => n24315);
   U17675 : INV_X1 port map( A => n24315, ZN => n24320);
   U17676 : MUX2_X1 port map( A => n24361, B => ADD_RD2(3), S => n22768, Z => 
                           n24319);
   U17677 : OAI21_X1 port map( B1 => n24320, B2 => CWP_3_port, A => n24319, ZN 
                           => n24314);
   U17678 : OAI21_X1 port map( B1 => n3043, B2 => n24315, A => n24314, ZN => 
                           n24318);
   U17679 : NOR2_X1 port map( A1 => n22768, A2 => n24360, ZN => n24316);
   U17680 : XOR2_X1 port map( A => n994, B => n24316, Z => n24317);
   U17681 : XOR2_X1 port map( A => n24318, B => n24317, Z => n16540);
   U17682 : XOR2_X1 port map( A => n24319, B => n3043, Z => n24321);
   U17683 : XOR2_X1 port map( A => n24321, B => n24320, Z => n25406);
   U17684 : INV_X1 port map( A => n25406, ZN => n16545);
   U17685 : NAND2_X1 port map( A1 => n24323, A2 => n24322, ZN => n24326);
   U17686 : INV_X1 port map( A => n24324, ZN => n24325);
   U17687 : XOR2_X1 port map( A => n24326, B => n24325, Z => n24335);
   U17688 : XOR2_X1 port map( A => n24327, B => n3046, Z => n24331);
   U17689 : INV_X1 port map( A => n24331, ZN => n24334);
   U17690 : XOR2_X1 port map( A => n24328, B => n3045, Z => n24330);
   U17691 : XOR2_X1 port map( A => n24330, B => n24329, Z => n24336);
   U17692 : INV_X1 port map( A => n24336, ZN => n24332);
   U17693 : INV_X1 port map( A => n24335, ZN => n24333);
   U17694 : OAI21_X1 port map( B1 => n3236, B2 => n23186, A => n24337, ZN => 
                           n5643);
   U17695 : OAI21_X1 port map( B1 => n3077, B2 => n24340, A => n24339, ZN => 
                           n5449);
   U17696 : NAND2_X1 port map( A1 => n24343, A2 => n23283, ZN => n25394);
   U17697 : NAND2_X1 port map( A1 => n22487, A2 => n22696, ZN => n24344);
   U17698 : NAND2_X1 port map( A1 => n22486, A2 => n22697, ZN => n24345);
   U17699 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), ZN => n24346
                           );
   U17700 : INV_X1 port map( A => n24346, ZN => n24352);
   U17701 : NAND2_X1 port map( A1 => n22696, A2 => ADD_RD1(0), ZN => n24347);
   U17702 : NAND2_X1 port map( A1 => n22697, A2 => n22484, ZN => n24376);
   U17703 : OAI222_X1 port map( A1 => n19676, A2 => n22516, B1 => n19548, B2 =>
                           n22935, C1 => n19612, C2 => n24376, ZN => n24348);
   U17704 : AOI221_X1 port map( B1 => n22970, B2 => n21284, C1 => n22912, C2 =>
                           n22225, A => n24348, ZN => n24375);
   U17705 : NAND3_X1 port map( A1 => n22484, A2 => n22696, A3 => n24369, ZN => 
                           n24349);
   U17706 : NAND3_X1 port map( A1 => n22696, A2 => n24369, A3 => n22486, ZN => 
                           n25388);
   U17707 : NAND3_X1 port map( A1 => N2739, A2 => n21456, A3 => n24350, ZN => 
                           n24351);
   U17708 : INV_X1 port map( A => n24351, ZN => n24356);
   U17709 : OAI22_X1 port map( A1 => n19228, A2 => n22965, B1 => n19164, B2 => 
                           n22976, ZN => n24353);
   U17710 : AOI221_X1 port map( B1 => n22803, B2 => n21286, C1 => n23268, C2 =>
                           n21841, A => n24353, ZN => n24374);
   U17711 : NAND3_X1 port map( A1 => n24356, A2 => n22484, A3 => n24369, ZN => 
                           n24354);
   U17712 : NAND3_X1 port map( A1 => n22932, A2 => ADD_RD1(2), A3 => n24368, ZN
                           => n25389);
   U17713 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => n22932
                           , ZN => n24386);
   U17714 : OAI222_X1 port map( A1 => n19100, A2 => n22635, B1 => n18972, B2 =>
                           n22951, C1 => n19036, C2 => n24386, ZN => n24357);
   U17715 : INV_X1 port map( A => n20769, ZN => n24358);
   U17716 : NAND2_X1 port map( A1 => n18513, A2 => n18514, ZN => n24363);
   U17717 : NAND2_X1 port map( A1 => n24361, A2 => n24360, ZN => n25371);
   U17718 : AOI21_X1 port map( B1 => n18517, B2 => n18518, A => n23196, ZN => 
                           n24362);
   U17719 : AOI221_X1 port map( B1 => n23212, B2 => n21907, C1 => n23204, C2 =>
                           n24363, A => n24362, ZN => n24367);
   U17720 : AOI222_X1 port map( A1 => n23236, A2 => n21350, B1 => n23228, B2 =>
                           n21026, C1 => n23220, C2 => n20833, ZN => n24366);
   U17721 : OAI222_X1 port map( A1 => n20444, A2 => n23260, B1 => n20572, B2 =>
                           n23252, C1 => n20508, C2 => n23244, ZN => n24364);
   U17722 : NOR4_X1 port map( A1 => n24364, A2 => n18523, A3 => n18509, A4 => 
                           n18510, ZN => n24365);
   U17723 : NAND3_X1 port map( A1 => n24367, A2 => n24366, A3 => n24365, ZN => 
                           n24371);
   U17724 : NAND3_X1 port map( A1 => n22488, A2 => n24369, A3 => n24368, ZN => 
                           n25392);
   U17725 : NAND3_X1 port map( A1 => n22488, A2 => ADD_RD1(0), A3 => n24369, ZN
                           => n24388);
   U17726 : OAI22_X1 port map( A1 => n18716, A2 => n22944, B1 => n18780, B2 => 
                           n24388, ZN => n24370);
   U17727 : AOI221_X1 port map( B1 => n22909, B2 => n24371, C1 => OUT1_0_port, 
                           C2 => n23271, A => n24370, ZN => n24372);
   U17728 : NAND4_X1 port map( A1 => n24375, A2 => n24374, A3 => n24373, A4 => 
                           n24372, ZN => n3275);
   U17729 : NAND2_X1 port map( A1 => n18474, A2 => n18475, ZN => n24378);
   U17730 : AOI21_X1 port map( B1 => n18478, B2 => n18479, A => n23196, ZN => 
                           n24377);
   U17731 : AOI221_X1 port map( B1 => n23212, B2 => n21844, C1 => n23204, C2 =>
                           n24378, A => n24377, ZN => n24382);
   U17732 : AOI222_X1 port map( A1 => n23236, A2 => n21287, B1 => n23228, B2 =>
                           n20963, C1 => n23220, C2 => n20770, ZN => n24381);
   U17733 : OAI222_X1 port map( A1 => n20443, A2 => n23260, B1 => n20571, B2 =>
                           n23252, C1 => n20507, C2 => n23244, ZN => n24379);
   U17734 : NOR4_X1 port map( A1 => n24379, A2 => n18483, A3 => n18470, A4 => 
                           n18471, ZN => n24380);
   U17735 : AND3_X1 port map( A1 => n24382, A2 => n24381, A3 => n24380, ZN => 
                           n24383);
   U17736 : OAI222_X1 port map( A1 => n19547, A2 => n22937, B1 => n24383, B2 =>
                           n22798, C1 => n19675, C2 => n22519, ZN => n24384);
   U17737 : AOI221_X1 port map( B1 => n22523, B2 => n22087, C1 => n22970, C2 =>
                           n21094, A => n24384, ZN => n24394);
   U17738 : OAI22_X1 port map( A1 => n19163, A2 => n22979, B1 => n19291, B2 => 
                           n22631, ZN => n24385);
   U17739 : AOI221_X1 port map( B1 => n22917, B2 => n22058, C1 => n22808, C2 =>
                           n21151, A => n24385, ZN => n24393);
   U17740 : OAI222_X1 port map( A1 => n18971, A2 => n22955, B1 => n19227, B2 =>
                           n22967, C1 => n19099, C2 => n22637, ZN => n24387);
   U17741 : AOI221_X1 port map( B1 => n25391, B2 => n22143, C1 => n22958, C2 =>
                           n21210, A => n24387, ZN => n24392);
   U17742 : OAI22_X1 port map( A1 => n23270, A2 => n24389, B1 => n18715, B2 => 
                           n22946, ZN => n24390);
   U17743 : AOI221_X1 port map( B1 => n23275, B2 => n20900, C1 => n22494, C2 =>
                           n21640, A => n24390, ZN => n24391);
   U17744 : NAND4_X1 port map( A1 => n24392, A2 => n24393, A3 => n24391, A4 => 
                           n24394, ZN => n3276);
   U17745 : NAND2_X1 port map( A1 => n18447, A2 => n18448, ZN => n24396);
   U17746 : AOI21_X1 port map( B1 => n18451, B2 => n18452, A => n23196, ZN => 
                           n24395);
   U17747 : AOI221_X1 port map( B1 => n23212, B2 => n21859, C1 => n23204, C2 =>
                           n24396, A => n24395, ZN => n24400);
   U17748 : AOI222_X1 port map( A1 => n23236, A2 => n21302, B1 => n23228, B2 =>
                           n20978, C1 => n23220, C2 => n20785, ZN => n24399);
   U17749 : OAI222_X1 port map( A1 => n20445, A2 => n23260, B1 => n20573, B2 =>
                           n23252, C1 => n20509, C2 => n23244, ZN => n24397);
   U17750 : NOR4_X1 port map( A1 => n24397, A2 => n18456, A3 => n18443, A4 => 
                           n18444, ZN => n24398);
   U17751 : AND3_X1 port map( A1 => n24400, A2 => n24399, A3 => n24398, ZN => 
                           n24401);
   U17752 : OAI222_X1 port map( A1 => n19549, A2 => n22936, B1 => n24401, B2 =>
                           n22800, C1 => n19677, C2 => n22517, ZN => n24402);
   U17753 : AOI221_X1 port map( B1 => n22921, B2 => n22088, C1 => n22971, C2 =>
                           n21109, A => n24402, ZN => n24410);
   U17754 : OAI22_X1 port map( A1 => n19165, A2 => n22978, B1 => n19293, B2 => 
                           n22648, ZN => n24403);
   U17755 : OAI222_X1 port map( A1 => n18973, A2 => n22954, B1 => n19229, B2 =>
                           n22965, C1 => n19101, C2 => n22636, ZN => n24404);
   U17756 : AOI221_X1 port map( B1 => n25391, B2 => n22037, C1 => n22959, C2 =>
                           n21225, A => n24404, ZN => n24408);
   U17757 : OAI22_X1 port map( A1 => n23270, A2 => n24405, B1 => n18717, B2 => 
                           n22947, ZN => n24406);
   U17758 : AOI221_X1 port map( B1 => n23275, B2 => n20914, C1 => n22494, C2 =>
                           n21654, A => n24406, ZN => n24407);
   U17759 : NAND4_X1 port map( A1 => n24407, A2 => n24409, A3 => n24408, A4 => 
                           n24410, ZN => n3277);
   U17760 : NAND2_X1 port map( A1 => n18420, A2 => n18421, ZN => n24412);
   U17761 : AOI21_X1 port map( B1 => n18424, B2 => n18425, A => n23196, ZN => 
                           n24411);
   U17762 : AOI221_X1 port map( B1 => n23212, B2 => n21860, C1 => n23204, C2 =>
                           n24412, A => n24411, ZN => n24416);
   U17763 : AOI222_X1 port map( A1 => n23236, A2 => n21303, B1 => n23228, B2 =>
                           n20979, C1 => n23220, C2 => n20786, ZN => n24415);
   U17764 : OAI222_X1 port map( A1 => n20442, A2 => n23260, B1 => n20570, B2 =>
                           n23252, C1 => n20506, C2 => n23244, ZN => n24413);
   U17765 : NOR4_X1 port map( A1 => n24413, A2 => n18429, A3 => n18416, A4 => 
                           n18417, ZN => n24414);
   U17766 : AND3_X1 port map( A1 => n24416, A2 => n24415, A3 => n24414, ZN => 
                           n24417);
   U17767 : OAI222_X1 port map( A1 => n19546, A2 => n22933, B1 => n24417, B2 =>
                           n22800, C1 => n19674, C2 => n22519, ZN => n24418);
   U17768 : AOI221_X1 port map( B1 => n22923, B2 => n22089, C1 => n22972, C2 =>
                           n21110, A => n24418, ZN => n24426);
   U17769 : OAI22_X1 port map( A1 => n19162, A2 => n22977, B1 => n19290, B2 => 
                           n22643, ZN => n24419);
   U17770 : AOI221_X1 port map( B1 => n22918, B2 => n22059, C1 => n22806, C2 =>
                           n21158, A => n24419, ZN => n24425);
   U17771 : OAI222_X1 port map( A1 => n18970, A2 => n22951, B1 => n19226, B2 =>
                           n22967, C1 => n19098, C2 => n22635, ZN => n24420);
   U17772 : AOI221_X1 port map( B1 => n22801, B2 => n22038, C1 => n22960, C2 =>
                           n21226, A => n24420, ZN => n24424);
   U17773 : OAI22_X1 port map( A1 => n23270, A2 => n24421, B1 => n18714, B2 => 
                           n22943, ZN => n24422);
   U17774 : AOI221_X1 port map( B1 => n23275, B2 => n20915, C1 => n22494, C2 =>
                           n21655, A => n24422, ZN => n24423);
   U17775 : NAND4_X1 port map( A1 => n24423, A2 => n24425, A3 => n24424, A4 => 
                           n24426, ZN => n3278);
   U17776 : NAND2_X1 port map( A1 => n18393, A2 => n18394, ZN => n24428);
   U17777 : AOI21_X1 port map( B1 => n18397, B2 => n18398, A => n23196, ZN => 
                           n24427);
   U17778 : AOI221_X1 port map( B1 => n23212, B2 => n21861, C1 => n23204, C2 =>
                           n24428, A => n24427, ZN => n24432);
   U17779 : AOI222_X1 port map( A1 => n23236, A2 => n21304, B1 => n23228, B2 =>
                           n20980, C1 => n23220, C2 => n20787, ZN => n24431);
   U17780 : OAI222_X1 port map( A1 => n20446, A2 => n23260, B1 => n20574, B2 =>
                           n23252, C1 => n20510, C2 => n23244, ZN => n24429);
   U17781 : NOR4_X1 port map( A1 => n24429, A2 => n18402, A3 => n18389, A4 => 
                           n18390, ZN => n24430);
   U17782 : AND3_X1 port map( A1 => n24432, A2 => n24431, A3 => n24430, ZN => 
                           n24433);
   U17783 : OAI222_X1 port map( A1 => n19550, A2 => n22936, B1 => n24433, B2 =>
                           n22800, C1 => n19678, C2 => n22516, ZN => n24434);
   U17784 : AOI221_X1 port map( B1 => n22923, B2 => n22090, C1 => n22971, C2 =>
                           n21111, A => n24434, ZN => n24442);
   U17785 : OAI22_X1 port map( A1 => n19166, A2 => n22976, B1 => n19294, B2 => 
                           n22634, ZN => n24435);
   U17786 : OAI222_X1 port map( A1 => n18974, A2 => n22953, B1 => n19230, B2 =>
                           n22966, C1 => n19102, C2 => n22639, ZN => n24436);
   U17787 : AOI221_X1 port map( B1 => n25391, B2 => n22144, C1 => n22962, C2 =>
                           n21227, A => n24436, ZN => n24440);
   U17788 : OAI22_X1 port map( A1 => n23270, A2 => n24437, B1 => n18718, B2 => 
                           n22943, ZN => n24438);
   U17789 : AOI221_X1 port map( B1 => n23275, B2 => n20916, C1 => n22494, C2 =>
                           n21656, A => n24438, ZN => n24439);
   U17790 : NAND4_X1 port map( A1 => n24440, A2 => n24441, A3 => n24439, A4 => 
                           n24442, ZN => n3279);
   U17791 : NAND2_X1 port map( A1 => n18366, A2 => n18367, ZN => n24444);
   U17792 : AOI21_X1 port map( B1 => n18370, B2 => n18371, A => n23196, ZN => 
                           n24443);
   U17793 : AOI221_X1 port map( B1 => n23212, B2 => n21845, C1 => n23204, C2 =>
                           n24444, A => n24443, ZN => n24448);
   U17794 : AOI222_X1 port map( A1 => n23236, A2 => n21288, B1 => n23228, B2 =>
                           n20964, C1 => n23220, C2 => n20771, ZN => n24447);
   U17795 : OAI222_X1 port map( A1 => n20441, A2 => n23260, B1 => n20569, B2 =>
                           n23252, C1 => n20505, C2 => n23244, ZN => n24445);
   U17796 : NOR4_X1 port map( A1 => n24445, A2 => n18375, A3 => n18362, A4 => 
                           n18363, ZN => n24446);
   U17797 : AND3_X1 port map( A1 => n24448, A2 => n24447, A3 => n24446, ZN => 
                           n24449);
   U17798 : OAI222_X1 port map( A1 => n19545, A2 => n22937, B1 => n24449, B2 =>
                           n22798, C1 => n19673, C2 => n22516, ZN => n24450);
   U17799 : AOI221_X1 port map( B1 => n22522, B2 => n22091, C1 => n22972, C2 =>
                           n21095, A => n24450, ZN => n24458);
   U17800 : OAI22_X1 port map( A1 => n19161, A2 => n22977, B1 => n19289, B2 => 
                           n22648, ZN => n24451);
   U17801 : OAI222_X1 port map( A1 => n18969, A2 => n22954, B1 => n19225, B2 =>
                           n22967, C1 => n19097, C2 => n22638, ZN => n24452);
   U17802 : AOI221_X1 port map( B1 => n25391, B2 => n22145, C1 => n22962, C2 =>
                           n21211, A => n24452, ZN => n24456);
   U17803 : OAI22_X1 port map( A1 => n23269, A2 => n24453, B1 => n18713, B2 => 
                           n22944, ZN => n24454);
   U17804 : AOI221_X1 port map( B1 => n23275, B2 => n20901, C1 => n22494, C2 =>
                           n21641, A => n24454, ZN => n24455);
   U17805 : NAND4_X1 port map( A1 => n24456, A2 => n24457, A3 => n24455, A4 => 
                           n24458, ZN => n3280);
   U17806 : NAND2_X1 port map( A1 => n18339, A2 => n18340, ZN => n24460);
   U17807 : AOI21_X1 port map( B1 => n18343, B2 => n18344, A => n23196, ZN => 
                           n24459);
   U17808 : AOI221_X1 port map( B1 => n23212, B2 => n21862, C1 => n23204, C2 =>
                           n24460, A => n24459, ZN => n24464);
   U17809 : AOI222_X1 port map( A1 => n23236, A2 => n21305, B1 => n23228, B2 =>
                           n20981, C1 => n23220, C2 => n20788, ZN => n24463);
   U17810 : OAI222_X1 port map( A1 => n20447, A2 => n23260, B1 => n20575, B2 =>
                           n23252, C1 => n20511, C2 => n23244, ZN => n24461);
   U17811 : NOR4_X1 port map( A1 => n24461, A2 => n18348, A3 => n18335, A4 => 
                           n18336, ZN => n24462);
   U17812 : AND3_X1 port map( A1 => n24464, A2 => n24463, A3 => n24462, ZN => 
                           n24465);
   U17813 : OAI222_X1 port map( A1 => n19551, A2 => n22933, B1 => n24465, B2 =>
                           n22800, C1 => n19679, C2 => n22517, ZN => n24466);
   U17814 : AOI221_X1 port map( B1 => n22522, B2 => n22092, C1 => n22973, C2 =>
                           n21112, A => n24466, ZN => n24474);
   U17815 : OAI22_X1 port map( A1 => n19167, A2 => n22978, B1 => n19295, B2 => 
                           n22647, ZN => n24467);
   U17816 : OAI222_X1 port map( A1 => n18975, A2 => n22954, B1 => n19231, B2 =>
                           n22964, C1 => n19103, C2 => n22638, ZN => n24468);
   U17817 : AOI221_X1 port map( B1 => n25391, B2 => n22146, C1 => n22962, C2 =>
                           n21228, A => n24468, ZN => n24472);
   U17818 : OAI22_X1 port map( A1 => n25394, A2 => n24469, B1 => n18719, B2 => 
                           n22945, ZN => n24470);
   U17819 : AOI221_X1 port map( B1 => n23275, B2 => n20917, C1 => n22494, C2 =>
                           n21657, A => n24470, ZN => n24471);
   U17820 : NAND4_X1 port map( A1 => n24472, A2 => n24473, A3 => n24471, A4 => 
                           n24474, ZN => n3281);
   U17821 : NAND2_X1 port map( A1 => n18312, A2 => n18313, ZN => n24476);
   U17822 : AOI21_X1 port map( B1 => n18316, B2 => n18317, A => n23196, ZN => 
                           n24475);
   U17823 : AOI221_X1 port map( B1 => n23212, B2 => n21877, C1 => n23204, C2 =>
                           n24476, A => n24475, ZN => n24480);
   U17824 : AOI222_X1 port map( A1 => n23236, A2 => n21320, B1 => n23228, B2 =>
                           n20996, C1 => n23220, C2 => n20803, ZN => n24479);
   U17825 : OAI222_X1 port map( A1 => n20440, A2 => n23260, B1 => n20568, B2 =>
                           n23252, C1 => n20504, C2 => n23244, ZN => n24477);
   U17826 : NOR4_X1 port map( A1 => n24477, A2 => n18321, A3 => n18308, A4 => 
                           n18309, ZN => n24478);
   U17827 : AND3_X1 port map( A1 => n24480, A2 => n24479, A3 => n24478, ZN => 
                           n24481);
   U17828 : OAI222_X1 port map( A1 => n19544, A2 => n22937, B1 => n24481, B2 =>
                           n22799, C1 => n19672, C2 => n22518, ZN => n24482);
   U17829 : AOI221_X1 port map( B1 => n22522, B2 => n22093, C1 => n22975, C2 =>
                           n21126, A => n24482, ZN => n24490);
   U17830 : OAI22_X1 port map( A1 => n19160, A2 => n22980, B1 => n19288, B2 => 
                           n22643, ZN => n24483);
   U17831 : AOI221_X1 port map( B1 => n22914, B2 => n22060, C1 => n22803, C2 =>
                           n21164, A => n24483, ZN => n24489);
   U17832 : OAI222_X1 port map( A1 => n18968, A2 => n22953, B1 => n19224, B2 =>
                           n22967, C1 => n19096, C2 => n22638, ZN => n24484);
   U17833 : AOI221_X1 port map( B1 => n25391, B2 => n22147, C1 => n22958, C2 =>
                           n21244, A => n24484, ZN => n24488);
   U17834 : OAI22_X1 port map( A1 => n23269, A2 => n24485, B1 => n18712, B2 => 
                           n22946, ZN => n24486);
   U17835 : AOI221_X1 port map( B1 => n23275, B2 => n20932, C1 => n22494, C2 =>
                           n21672, A => n24486, ZN => n24487);
   U17836 : NAND4_X1 port map( A1 => n24488, A2 => n24489, A3 => n24487, A4 => 
                           n24490, ZN => n3282);
   U17837 : NAND2_X1 port map( A1 => n18285, A2 => n18286, ZN => n24492);
   U17838 : AOI21_X1 port map( B1 => n18289, B2 => n18290, A => n23196, ZN => 
                           n24491);
   U17839 : AOI221_X1 port map( B1 => n23212, B2 => n21878, C1 => n23204, C2 =>
                           n24492, A => n24491, ZN => n24496);
   U17840 : AOI222_X1 port map( A1 => n23236, A2 => n21321, B1 => n23228, B2 =>
                           n20997, C1 => n23220, C2 => n20804, ZN => n24495);
   U17841 : OAI222_X1 port map( A1 => n20448, A2 => n23260, B1 => n20576, B2 =>
                           n23252, C1 => n20512, C2 => n23244, ZN => n24493);
   U17842 : NOR4_X1 port map( A1 => n24493, A2 => n18294, A3 => n18281, A4 => 
                           n18282, ZN => n24494);
   U17843 : AND3_X1 port map( A1 => n24496, A2 => n24495, A3 => n24494, ZN => 
                           n24497);
   U17844 : OAI222_X1 port map( A1 => n19552, A2 => n22935, B1 => n24497, B2 =>
                           n22799, C1 => n19680, C2 => n22518, ZN => n24498);
   U17845 : AOI221_X1 port map( B1 => n22923, B2 => n22094, C1 => n22970, C2 =>
                           n21127, A => n24498, ZN => n24506);
   U17846 : OAI22_X1 port map( A1 => n19168, A2 => n22979, B1 => n19296, B2 => 
                           n22647, ZN => n24499);
   U17847 : OAI222_X1 port map( A1 => n18976, A2 => n22953, B1 => n19232, B2 =>
                           n22964, C1 => n19104, C2 => n22639, ZN => n24500);
   U17848 : AOI221_X1 port map( B1 => n25391, B2 => n22148, C1 => n22959, C2 =>
                           n21245, A => n24500, ZN => n24504);
   U17849 : OAI22_X1 port map( A1 => n25394, A2 => n24501, B1 => n18720, B2 => 
                           n22945, ZN => n24502);
   U17850 : AOI221_X1 port map( B1 => n23275, B2 => n20933, C1 => n22494, C2 =>
                           n21673, A => n24502, ZN => n24503);
   U17851 : NAND4_X1 port map( A1 => n24504, A2 => n24505, A3 => n24503, A4 => 
                           n24506, ZN => n3283);
   U17852 : NAND2_X1 port map( A1 => n18258, A2 => n18259, ZN => n24508);
   U17853 : AOI21_X1 port map( B1 => n18262, B2 => n18263, A => n23196, ZN => 
                           n24507);
   U17854 : AOI221_X1 port map( B1 => n23212, B2 => n21900, C1 => n23204, C2 =>
                           n24508, A => n24507, ZN => n24512);
   U17855 : AOI222_X1 port map( A1 => n23236, A2 => n21343, B1 => n23228, B2 =>
                           n21019, C1 => n23220, C2 => n20826, ZN => n24511);
   U17856 : OAI222_X1 port map( A1 => n20439, A2 => n23260, B1 => n20567, B2 =>
                           n23252, C1 => n20503, C2 => n23244, ZN => n24509);
   U17857 : NOR4_X1 port map( A1 => n24509, A2 => n18267, A3 => n18254, A4 => 
                           n18255, ZN => n24510);
   U17858 : AND3_X1 port map( A1 => n24512, A2 => n24511, A3 => n24510, ZN => 
                           n24513);
   U17859 : OAI222_X1 port map( A1 => n19543, A2 => n22652, B1 => n24513, B2 =>
                           n22799, C1 => n19671, C2 => n22519, ZN => n24514);
   U17860 : AOI221_X1 port map( B1 => n22923, B2 => n22184, C1 => n22971, C2 =>
                           n21150, A => n24514, ZN => n24522);
   U17861 : OAI22_X1 port map( A1 => n19159, A2 => n22978, B1 => n19287, B2 => 
                           n22651, ZN => n24515);
   U17862 : OAI222_X1 port map( A1 => n18967, A2 => n22952, B1 => n19223, B2 =>
                           n22966, C1 => n19095, C2 => n22635, ZN => n24516);
   U17863 : AOI221_X1 port map( B1 => n22801, B2 => n22039, C1 => n22957, C2 =>
                           n21266, A => n24516, ZN => n24520);
   U17864 : OAI22_X1 port map( A1 => n25394, A2 => n24517, B1 => n18711, B2 => 
                           n22946, ZN => n24518);
   U17865 : AOI221_X1 port map( B1 => n23275, B2 => n20955, C1 => n22494, C2 =>
                           n21751, A => n24518, ZN => n24519);
   U17866 : NAND4_X1 port map( A1 => n24522, A2 => n24521, A3 => n24520, A4 => 
                           n24519, ZN => n3284);
   U17867 : NAND2_X1 port map( A1 => n18231, A2 => n18232, ZN => n24524);
   U17868 : AOI21_X1 port map( B1 => n18235, B2 => n18236, A => n23196, ZN => 
                           n24523);
   U17869 : AOI221_X1 port map( B1 => n23212, B2 => n21879, C1 => n23204, C2 =>
                           n24524, A => n24523, ZN => n24528);
   U17870 : AOI222_X1 port map( A1 => n23236, A2 => n21322, B1 => n23228, B2 =>
                           n20998, C1 => n23220, C2 => n20805, ZN => n24527);
   U17871 : OAI222_X1 port map( A1 => n20449, A2 => n23260, B1 => n20577, B2 =>
                           n23252, C1 => n20513, C2 => n23244, ZN => n24525);
   U17872 : NOR4_X1 port map( A1 => n24525, A2 => n18240, A3 => n18227, A4 => 
                           n18228, ZN => n24526);
   U17873 : AND3_X1 port map( A1 => n24528, A2 => n24527, A3 => n24526, ZN => 
                           n24529);
   U17874 : OAI222_X1 port map( A1 => n19553, A2 => n22933, B1 => n24529, B2 =>
                           n22799, C1 => n19681, C2 => n22521, ZN => n24530);
   U17875 : AOI221_X1 port map( B1 => n22522, B2 => n22095, C1 => n22972, C2 =>
                           n21128, A => n24530, ZN => n24538);
   U17876 : OAI22_X1 port map( A1 => n19169, A2 => n22976, B1 => n19297, B2 => 
                           n22631, ZN => n24531);
   U17877 : AOI221_X1 port map( B1 => n22920, B2 => n22061, C1 => n22802, C2 =>
                           n21165, A => n24531, ZN => n24537);
   U17878 : OAI222_X1 port map( A1 => n18977, A2 => n22955, B1 => n19233, B2 =>
                           n22964, C1 => n19105, C2 => n22637, ZN => n24532);
   U17879 : AOI221_X1 port map( B1 => n25391, B2 => n22149, C1 => n22958, C2 =>
                           n21246, A => n24532, ZN => n24536);
   U17880 : OAI22_X1 port map( A1 => n23269, A2 => n24533, B1 => n18721, B2 => 
                           n22947, ZN => n24534);
   U17881 : AOI221_X1 port map( B1 => n23275, B2 => n20934, C1 => n22494, C2 =>
                           n21674, A => n24534, ZN => n24535);
   U17882 : NAND4_X1 port map( A1 => n24536, A2 => n24537, A3 => n24535, A4 => 
                           n24538, ZN => n3285);
   U17883 : NAND2_X1 port map( A1 => n18204, A2 => n18205, ZN => n24540);
   U17884 : AOI21_X1 port map( B1 => n18208, B2 => n18209, A => n23196, ZN => 
                           n24539);
   U17885 : AOI221_X1 port map( B1 => n23212, B2 => n21863, C1 => n23204, C2 =>
                           n24540, A => n24539, ZN => n24544);
   U17886 : AOI222_X1 port map( A1 => n23236, A2 => n21306, B1 => n23228, B2 =>
                           n20982, C1 => n23220, C2 => n20789, ZN => n24543);
   U17887 : OAI222_X1 port map( A1 => n20438, A2 => n23260, B1 => n20566, B2 =>
                           n23252, C1 => n20502, C2 => n23244, ZN => n24541);
   U17888 : NOR4_X1 port map( A1 => n24541, A2 => n18213, A3 => n18200, A4 => 
                           n18201, ZN => n24542);
   U17889 : AND3_X1 port map( A1 => n24544, A2 => n24543, A3 => n24542, ZN => 
                           n24545);
   U17890 : OAI222_X1 port map( A1 => n19542, A2 => n22936, B1 => n24545, B2 =>
                           n22800, C1 => n19670, C2 => n22520, ZN => n24546);
   U17891 : AOI221_X1 port map( B1 => n22523, B2 => n22096, C1 => n22973, C2 =>
                           n21113, A => n24546, ZN => n24554);
   U17892 : OAI22_X1 port map( A1 => n19158, A2 => n22977, B1 => n19286, B2 => 
                           n22634, ZN => n24547);
   U17893 : AOI221_X1 port map( B1 => n22917, B2 => n22062, C1 => n22811, C2 =>
                           n21159, A => n24547, ZN => n24553);
   U17894 : OAI222_X1 port map( A1 => n18966, A2 => n22952, B1 => n19222, B2 =>
                           n22968, C1 => n19094, C2 => n22635, ZN => n24548);
   U17895 : AOI221_X1 port map( B1 => n25391, B2 => n22150, C1 => n22959, C2 =>
                           n21229, A => n24548, ZN => n24552);
   U17896 : OAI22_X1 port map( A1 => n23270, A2 => n24549, B1 => n18710, B2 => 
                           n22943, ZN => n24550);
   U17897 : AOI221_X1 port map( B1 => n23275, B2 => n20918, C1 => n22494, C2 =>
                           n21658, A => n24550, ZN => n24551);
   U17898 : NAND4_X1 port map( A1 => n24552, A2 => n24553, A3 => n24551, A4 => 
                           n24554, ZN => n3286);
   U17899 : NAND2_X1 port map( A1 => n18177, A2 => n18178, ZN => n24556);
   U17900 : AOI21_X1 port map( B1 => n18181, B2 => n18182, A => n23197, ZN => 
                           n24555);
   U17901 : AOI221_X1 port map( B1 => n23213, B2 => n21864, C1 => n23205, C2 =>
                           n24556, A => n24555, ZN => n24560);
   U17902 : AOI222_X1 port map( A1 => n23237, A2 => n21307, B1 => n23229, B2 =>
                           n20983, C1 => n23221, C2 => n20790, ZN => n24559);
   U17903 : OAI222_X1 port map( A1 => n20450, A2 => n23261, B1 => n20578, B2 =>
                           n23253, C1 => n20514, C2 => n23245, ZN => n24557);
   U17904 : NOR4_X1 port map( A1 => n24557, A2 => n18186, A3 => n18173, A4 => 
                           n18174, ZN => n24558);
   U17905 : AND3_X1 port map( A1 => n24560, A2 => n24559, A3 => n24558, ZN => 
                           n24561);
   U17906 : OAI222_X1 port map( A1 => n19554, A2 => n22937, B1 => n24561, B2 =>
                           n22800, C1 => n19682, C2 => n22517, ZN => n24562);
   U17907 : AOI221_X1 port map( B1 => n22523, B2 => n22097, C1 => n22974, C2 =>
                           n21114, A => n24562, ZN => n24570);
   U17908 : OAI22_X1 port map( A1 => n19170, A2 => n22977, B1 => n19298, B2 => 
                           n22650, ZN => n24563);
   U17909 : OAI222_X1 port map( A1 => n18978, A2 => n22955, B1 => n19234, B2 =>
                           n22967, C1 => n19106, C2 => n22638, ZN => n24564);
   U17910 : AOI221_X1 port map( B1 => n25391, B2 => n22151, C1 => n22960, C2 =>
                           n21230, A => n24564, ZN => n24568);
   U17911 : OAI22_X1 port map( A1 => n23270, A2 => n24565, B1 => n18722, B2 => 
                           n22947, ZN => n24566);
   U17912 : AOI221_X1 port map( B1 => n23276, B2 => n20919, C1 => n22494, C2 =>
                           n21659, A => n24566, ZN => n24567);
   U17913 : NAND4_X1 port map( A1 => n24568, A2 => n24569, A3 => n24567, A4 => 
                           n24570, ZN => n3287);
   U17914 : NAND2_X1 port map( A1 => n18150, A2 => n18151, ZN => n24572);
   U17915 : AOI21_X1 port map( B1 => n18154, B2 => n18155, A => n23197, ZN => 
                           n24571);
   U17916 : AOI221_X1 port map( B1 => n23213, B2 => n21880, C1 => n23205, C2 =>
                           n24572, A => n24571, ZN => n24576);
   U17917 : AOI222_X1 port map( A1 => n23237, A2 => n21323, B1 => n23229, B2 =>
                           n20999, C1 => n23221, C2 => n20806, ZN => n24575);
   U17918 : OAI222_X1 port map( A1 => n20437, A2 => n23261, B1 => n20565, B2 =>
                           n23253, C1 => n20501, C2 => n23245, ZN => n24573);
   U17919 : NOR4_X1 port map( A1 => n24573, A2 => n18159, A3 => n18146, A4 => 
                           n18147, ZN => n24574);
   U17920 : AND3_X1 port map( A1 => n24576, A2 => n24575, A3 => n24574, ZN => 
                           n24577);
   U17921 : OAI222_X1 port map( A1 => n19541, A2 => n22937, B1 => n24577, B2 =>
                           n22799, C1 => n19669, C2 => n22520, ZN => n24578);
   U17922 : AOI221_X1 port map( B1 => n22921, B2 => n22098, C1 => n22970, C2 =>
                           n21129, A => n24578, ZN => n24586);
   U17923 : OAI22_X1 port map( A1 => n19157, A2 => n22976, B1 => n19285, B2 => 
                           n22651, ZN => n24579);
   U17924 : OAI222_X1 port map( A1 => n18965, A2 => n22955, B1 => n19221, B2 =>
                           n22968, C1 => n19093, C2 => n22639, ZN => n24580);
   U17925 : AOI221_X1 port map( B1 => n25391, B2 => n22152, C1 => n22961, C2 =>
                           n21247, A => n24580, ZN => n24584);
   U17926 : OAI22_X1 port map( A1 => n25394, A2 => n24581, B1 => n18709, B2 => 
                           n22946, ZN => n24582);
   U17927 : AOI221_X1 port map( B1 => n23276, B2 => n20935, C1 => n22494, C2 =>
                           n21675, A => n24582, ZN => n24583);
   U17928 : NAND4_X1 port map( A1 => n24584, A2 => n24585, A3 => n24583, A4 => 
                           n24586, ZN => n3288);
   U17929 : NAND2_X1 port map( A1 => n18123, A2 => n18124, ZN => n24588);
   U17930 : AOI21_X1 port map( B1 => n18127, B2 => n18128, A => n23197, ZN => 
                           n24587);
   U17931 : AOI221_X1 port map( B1 => n23213, B2 => n21865, C1 => n23205, C2 =>
                           n24588, A => n24587, ZN => n24592);
   U17932 : AOI222_X1 port map( A1 => n23237, A2 => n21308, B1 => n23229, B2 =>
                           n20984, C1 => n23221, C2 => n20791, ZN => n24591);
   U17933 : OAI222_X1 port map( A1 => n20451, A2 => n23261, B1 => n20579, B2 =>
                           n23253, C1 => n20515, C2 => n23245, ZN => n24589);
   U17934 : NOR4_X1 port map( A1 => n24589, A2 => n18132, A3 => n18119, A4 => 
                           n18120, ZN => n24590);
   U17935 : AND3_X1 port map( A1 => n24592, A2 => n24591, A3 => n24590, ZN => 
                           n24593);
   U17936 : OAI222_X1 port map( A1 => n19555, A2 => n22935, B1 => n24593, B2 =>
                           n22800, C1 => n19683, C2 => n22519, ZN => n24594);
   U17937 : AOI221_X1 port map( B1 => n22923, B2 => n22099, C1 => n22974, C2 =>
                           n21115, A => n24594, ZN => n24602);
   U17938 : OAI22_X1 port map( A1 => n19171, A2 => n22980, B1 => n19299, B2 => 
                           n22641, ZN => n24595);
   U17939 : OAI222_X1 port map( A1 => n18979, A2 => n22953, B1 => n19235, B2 =>
                           n22968, C1 => n19107, C2 => n22638, ZN => n24596);
   U17940 : AOI221_X1 port map( B1 => n25391, B2 => n22153, C1 => n22962, C2 =>
                           n21231, A => n24596, ZN => n24600);
   U17941 : OAI22_X1 port map( A1 => n25394, A2 => n24597, B1 => n18723, B2 => 
                           n22944, ZN => n24598);
   U17942 : AOI221_X1 port map( B1 => n23276, B2 => n20920, C1 => n22494, C2 =>
                           n21660, A => n24598, ZN => n24599);
   U17943 : NAND4_X1 port map( A1 => n24600, A2 => n24601, A3 => n24599, A4 => 
                           n24602, ZN => n3289);
   U17944 : NAND2_X1 port map( A1 => n18096, A2 => n18097, ZN => n24604);
   U17945 : AOI21_X1 port map( B1 => n18100, B2 => n18101, A => n23197, ZN => 
                           n24603);
   U17946 : AOI221_X1 port map( B1 => n23213, B2 => n21902, C1 => n23205, C2 =>
                           n24604, A => n24603, ZN => n24608);
   U17947 : AOI222_X1 port map( A1 => n23237, A2 => n21345, B1 => n23229, B2 =>
                           n21021, C1 => n23221, C2 => n20828, ZN => n24607);
   U17948 : OAI222_X1 port map( A1 => n20436, A2 => n23261, B1 => n20564, B2 =>
                           n23253, C1 => n20500, C2 => n23245, ZN => n24605);
   U17949 : NOR4_X1 port map( A1 => n24605, A2 => n18105, A3 => n18092, A4 => 
                           n18093, ZN => n24606);
   U17950 : AND3_X1 port map( A1 => n24608, A2 => n24607, A3 => n24606, ZN => 
                           n24609);
   U17951 : OAI222_X1 port map( A1 => n19540, A2 => n22933, B1 => n24609, B2 =>
                           n22798, C1 => n19668, C2 => n22517, ZN => n24610);
   U17952 : OAI22_X1 port map( A1 => n19156, A2 => n22980, B1 => n19284, B2 => 
                           n22644, ZN => n24611);
   U17953 : OAI222_X1 port map( A1 => n18964, A2 => n22951, B1 => n19220, B2 =>
                           n22966, C1 => n19092, C2 => n22635, ZN => n24612);
   U17954 : AOI221_X1 port map( B1 => n22801, B2 => n22040, C1 => n22962, C2 =>
                           n21279, A => n24612, ZN => n24616);
   U17955 : OAI22_X1 port map( A1 => n25394, A2 => n24613, B1 => n18708, B2 => 
                           n22945, ZN => n24614);
   U17956 : AOI221_X1 port map( B1 => n23276, B2 => n20957, C1 => n22494, C2 =>
                           n21830, A => n24614, ZN => n24615);
   U17957 : NAND4_X1 port map( A1 => n24615, A2 => n24617, A3 => n24616, A4 => 
                           n24618, ZN => n3290);
   U17958 : NAND2_X1 port map( A1 => n18069, A2 => n18070, ZN => n24620);
   U17959 : AOI21_X1 port map( B1 => n18073, B2 => n18074, A => n23197, ZN => 
                           n24619);
   U17960 : AOI221_X1 port map( B1 => n23213, B2 => n21866, C1 => n23205, C2 =>
                           n24620, A => n24619, ZN => n24624);
   U17961 : AOI222_X1 port map( A1 => n23237, A2 => n21309, B1 => n23229, B2 =>
                           n20985, C1 => n23221, C2 => n20792, ZN => n24623);
   U17962 : OAI222_X1 port map( A1 => n20452, A2 => n23261, B1 => n20580, B2 =>
                           n23253, C1 => n20516, C2 => n23245, ZN => n24621);
   U17963 : NOR4_X1 port map( A1 => n24621, A2 => n18078, A3 => n18065, A4 => 
                           n18066, ZN => n24622);
   U17964 : AND3_X1 port map( A1 => n24624, A2 => n24623, A3 => n24622, ZN => 
                           n24625);
   U17965 : OAI222_X1 port map( A1 => n19556, A2 => n22936, B1 => n24625, B2 =>
                           n22800, C1 => n19684, C2 => n22521, ZN => n24626);
   U17966 : AOI221_X1 port map( B1 => n22523, B2 => n22100, C1 => n22973, C2 =>
                           n21116, A => n24626, ZN => n24634);
   U17967 : OAI22_X1 port map( A1 => n19172, A2 => n22976, B1 => n19300, B2 => 
                           n22641, ZN => n24627);
   U17968 : OAI222_X1 port map( A1 => n18980, A2 => n22954, B1 => n19236, B2 =>
                           n22965, C1 => n19108, C2 => n22635, ZN => n24628);
   U17969 : AOI221_X1 port map( B1 => n25391, B2 => n22154, C1 => n22958, C2 =>
                           n21232, A => n24628, ZN => n24632);
   U17970 : OAI22_X1 port map( A1 => n23269, A2 => n24629, B1 => n18724, B2 => 
                           n22943, ZN => n24630);
   U17971 : AOI221_X1 port map( B1 => n23276, B2 => n20921, C1 => n22494, C2 =>
                           n21661, A => n24630, ZN => n24631);
   U17972 : NAND4_X1 port map( A1 => n24632, A2 => n24633, A3 => n24631, A4 => 
                           n24634, ZN => n3291);
   U17973 : NAND2_X1 port map( A1 => n18042, A2 => n18043, ZN => n24636);
   U17974 : AOI21_X1 port map( B1 => n18046, B2 => n18047, A => n23197, ZN => 
                           n24635);
   U17975 : AOI221_X1 port map( B1 => n23213, B2 => n21881, C1 => n23205, C2 =>
                           n24636, A => n24635, ZN => n24640);
   U17976 : AOI222_X1 port map( A1 => n23237, A2 => n21324, B1 => n23229, B2 =>
                           n21000, C1 => n23221, C2 => n20807, ZN => n24639);
   U17977 : OAI222_X1 port map( A1 => n20435, A2 => n23261, B1 => n20563, B2 =>
                           n23253, C1 => n20499, C2 => n23245, ZN => n24637);
   U17978 : NOR4_X1 port map( A1 => n24637, A2 => n18051, A3 => n18038, A4 => 
                           n18039, ZN => n24638);
   U17979 : AND3_X1 port map( A1 => n24640, A2 => n24639, A3 => n24638, ZN => 
                           n24641);
   U17980 : OAI222_X1 port map( A1 => n19539, A2 => n22652, B1 => n24641, B2 =>
                           n22799, C1 => n19667, C2 => n22519, ZN => n24642);
   U17981 : AOI221_X1 port map( B1 => n22522, B2 => n22101, C1 => n22974, C2 =>
                           n21130, A => n24642, ZN => n24650);
   U17982 : OAI22_X1 port map( A1 => n19155, A2 => n22979, B1 => n19283, B2 => 
                           n22634, ZN => n24643);
   U17983 : AOI221_X1 port map( B1 => n22917, B2 => n22063, C1 => n22807, C2 =>
                           n21166, A => n24643, ZN => n24649);
   U17984 : OAI222_X1 port map( A1 => n18963, A2 => n22954, B1 => n19219, B2 =>
                           n22965, C1 => n19091, C2 => n22637, ZN => n24644);
   U17985 : AOI221_X1 port map( B1 => n25391, B2 => n22155, C1 => n22957, C2 =>
                           n21248, A => n24644, ZN => n24648);
   U17986 : OAI22_X1 port map( A1 => n25394, A2 => n24645, B1 => n18707, B2 => 
                           n22946, ZN => n24646);
   U17987 : AOI221_X1 port map( B1 => n23276, B2 => n20936, C1 => n22494, C2 =>
                           n21676, A => n24646, ZN => n24647);
   U17988 : NAND4_X1 port map( A1 => n24648, A2 => n24649, A3 => n24647, A4 => 
                           n24650, ZN => n3292);
   U17989 : NAND2_X1 port map( A1 => n18015, A2 => n18016, ZN => n24652);
   U17990 : AOI21_X1 port map( B1 => n18019, B2 => n18020, A => n23197, ZN => 
                           n24651);
   U17991 : AOI221_X1 port map( B1 => n23213, B2 => n21867, C1 => n23205, C2 =>
                           n24652, A => n24651, ZN => n24656);
   U17992 : AOI222_X1 port map( A1 => n23237, A2 => n21310, B1 => n23229, B2 =>
                           n20986, C1 => n23221, C2 => n20793, ZN => n24655);
   U17993 : OAI222_X1 port map( A1 => n20453, A2 => n23261, B1 => n20581, B2 =>
                           n23253, C1 => n20517, C2 => n23245, ZN => n24653);
   U17994 : NOR4_X1 port map( A1 => n24653, A2 => n18024, A3 => n18011, A4 => 
                           n18012, ZN => n24654);
   U17995 : AND3_X1 port map( A1 => n24656, A2 => n24655, A3 => n24654, ZN => 
                           n24657);
   U17996 : OAI222_X1 port map( A1 => n19557, A2 => n22933, B1 => n24657, B2 =>
                           n22800, C1 => n19685, C2 => n22519, ZN => n24658);
   U17997 : AOI221_X1 port map( B1 => n22523, B2 => n22102, C1 => n22974, C2 =>
                           n21117, A => n24658, ZN => n24666);
   U17998 : OAI22_X1 port map( A1 => n19173, A2 => n22978, B1 => n19301, B2 => 
                           n22640, ZN => n24659);
   U17999 : AOI221_X1 port map( B1 => n22912, B2 => n22064, C1 => n22802, C2 =>
                           n21160, A => n24659, ZN => n24665);
   U18000 : OAI222_X1 port map( A1 => n18981, A2 => n22955, B1 => n19237, B2 =>
                           n22965, C1 => n19109, C2 => n22637, ZN => n24660);
   U18001 : AOI221_X1 port map( B1 => n22801, B2 => n22041, C1 => n22960, C2 =>
                           n21233, A => n24660, ZN => n24664);
   U18002 : OAI22_X1 port map( A1 => n23269, A2 => n24661, B1 => n18725, B2 => 
                           n22947, ZN => n24662);
   U18003 : AOI221_X1 port map( B1 => n23276, B2 => n20922, C1 => n22494, C2 =>
                           n21662, A => n24662, ZN => n24663);
   U18004 : NAND4_X1 port map( A1 => n24663, A2 => n24665, A3 => n24664, A4 => 
                           n24666, ZN => n3293);
   U18005 : NAND2_X1 port map( A1 => n17988, A2 => n17989, ZN => n24668);
   U18006 : AOI21_X1 port map( B1 => n17992, B2 => n17993, A => n23197, ZN => 
                           n24667);
   U18007 : AOI221_X1 port map( B1 => n23213, B2 => n21846, C1 => n23205, C2 =>
                           n24668, A => n24667, ZN => n24672);
   U18008 : AOI222_X1 port map( A1 => n23237, A2 => n21289, B1 => n23229, B2 =>
                           n20965, C1 => n23221, C2 => n20772, ZN => n24671);
   U18009 : OAI222_X1 port map( A1 => n20434, A2 => n23261, B1 => n20562, B2 =>
                           n23253, C1 => n20498, C2 => n23245, ZN => n24669);
   U18010 : NOR4_X1 port map( A1 => n24669, A2 => n17997, A3 => n17984, A4 => 
                           n17985, ZN => n24670);
   U18011 : AND3_X1 port map( A1 => n24672, A2 => n24671, A3 => n24670, ZN => 
                           n24673);
   U18012 : OAI222_X1 port map( A1 => n19538, A2 => n22935, B1 => n24673, B2 =>
                           n22798, C1 => n19666, C2 => n22518, ZN => n24674);
   U18013 : AOI221_X1 port map( B1 => n22922, B2 => n22103, C1 => n22972, C2 =>
                           n21096, A => n24674, ZN => n24682);
   U18014 : OAI22_X1 port map( A1 => n19154, A2 => n22977, B1 => n19282, B2 => 
                           n22649, ZN => n24675);
   U18015 : AOI221_X1 port map( B1 => n22912, B2 => n22065, C1 => n22809, C2 =>
                           n21152, A => n24675, ZN => n24681);
   U18016 : OAI222_X1 port map( A1 => n18962, A2 => n22953, B1 => n19218, B2 =>
                           n22964, C1 => n19090, C2 => n22635, ZN => n24676);
   U18017 : AOI221_X1 port map( B1 => n25391, B2 => n22156, C1 => n22962, C2 =>
                           n21212, A => n24676, ZN => n24680);
   U18018 : OAI22_X1 port map( A1 => n25394, A2 => n24677, B1 => n18706, B2 => 
                           n22944, ZN => n24678);
   U18019 : AOI221_X1 port map( B1 => n23276, B2 => n20902, C1 => n22494, C2 =>
                           n21642, A => n24678, ZN => n24679);
   U18020 : NAND4_X1 port map( A1 => n24680, A2 => n24681, A3 => n24679, A4 => 
                           n24682, ZN => n3294);
   U18021 : NAND2_X1 port map( A1 => n17961, A2 => n17962, ZN => n24684);
   U18022 : AOI21_X1 port map( B1 => n17965, B2 => n17966, A => n23197, ZN => 
                           n24683);
   U18023 : AOI221_X1 port map( B1 => n23213, B2 => n21868, C1 => n23205, C2 =>
                           n24684, A => n24683, ZN => n24688);
   U18024 : AOI222_X1 port map( A1 => n23237, A2 => n21311, B1 => n23229, B2 =>
                           n20987, C1 => n23221, C2 => n20794, ZN => n24687);
   U18025 : OAI222_X1 port map( A1 => n20454, A2 => n23261, B1 => n20582, B2 =>
                           n23253, C1 => n20518, C2 => n23245, ZN => n24685);
   U18026 : NOR4_X1 port map( A1 => n24685, A2 => n17970, A3 => n17957, A4 => 
                           n17958, ZN => n24686);
   U18027 : AND3_X1 port map( A1 => n24688, A2 => n24687, A3 => n24686, ZN => 
                           n24689);
   U18028 : OAI222_X1 port map( A1 => n19558, A2 => n22934, B1 => n24689, B2 =>
                           n22800, C1 => n19686, C2 => n22521, ZN => n24690);
   U18029 : AOI221_X1 port map( B1 => n22922, B2 => n22104, C1 => n22973, C2 =>
                           n21118, A => n24690, ZN => n24698);
   U18030 : OAI22_X1 port map( A1 => n19174, A2 => n22979, B1 => n19302, B2 => 
                           n22644, ZN => n24691);
   U18031 : OAI222_X1 port map( A1 => n18982, A2 => n22952, B1 => n19238, B2 =>
                           n22965, C1 => n19110, C2 => n22636, ZN => n24692);
   U18032 : AOI221_X1 port map( B1 => n25391, B2 => n22157, C1 => n22957, C2 =>
                           n21234, A => n24692, ZN => n24696);
   U18033 : OAI22_X1 port map( A1 => n23269, A2 => n24693, B1 => n18726, B2 => 
                           n22945, ZN => n24694);
   U18034 : AOI221_X1 port map( B1 => n23276, B2 => n20923, C1 => n22494, C2 =>
                           n21663, A => n24694, ZN => n24695);
   U18035 : NAND4_X1 port map( A1 => n24696, A2 => n24697, A3 => n24695, A4 => 
                           n24698, ZN => n3295);
   U18036 : NAND2_X1 port map( A1 => n17934, A2 => n17935, ZN => n24700);
   U18037 : AOI21_X1 port map( B1 => n17938, B2 => n17939, A => n23197, ZN => 
                           n24699);
   U18038 : AOI221_X1 port map( B1 => n23213, B2 => n21882, C1 => n23205, C2 =>
                           n24700, A => n24699, ZN => n24704);
   U18039 : AOI222_X1 port map( A1 => n23237, A2 => n21325, B1 => n23229, B2 =>
                           n21001, C1 => n23221, C2 => n20808, ZN => n24703);
   U18040 : OAI222_X1 port map( A1 => n20433, A2 => n23261, B1 => n20561, B2 =>
                           n23253, C1 => n20497, C2 => n23245, ZN => n24701);
   U18041 : NOR4_X1 port map( A1 => n24701, A2 => n17943, A3 => n17930, A4 => 
                           n17931, ZN => n24702);
   U18042 : AND3_X1 port map( A1 => n24704, A2 => n24703, A3 => n24702, ZN => 
                           n24705);
   U18043 : OAI222_X1 port map( A1 => n19537, A2 => n22937, B1 => n24705, B2 =>
                           n22799, C1 => n19665, C2 => n22520, ZN => n24706);
   U18044 : AOI221_X1 port map( B1 => n22921, B2 => n22105, C1 => n22974, C2 =>
                           n21131, A => n24706, ZN => n24714);
   U18045 : OAI22_X1 port map( A1 => n19153, A2 => n22980, B1 => n19281, B2 => 
                           n22640, ZN => n24707);
   U18046 : AOI221_X1 port map( B1 => n22913, B2 => n22066, C1 => n22811, C2 =>
                           n21167, A => n24707, ZN => n24713);
   U18047 : OAI222_X1 port map( A1 => n18961, A2 => n22952, B1 => n19217, B2 =>
                           n22968, C1 => n19089, C2 => n22639, ZN => n24708);
   U18048 : AOI221_X1 port map( B1 => n25391, B2 => n22158, C1 => n22962, C2 =>
                           n21249, A => n24708, ZN => n24712);
   U18049 : OAI22_X1 port map( A1 => n25394, A2 => n24709, B1 => n18705, B2 => 
                           n22946, ZN => n24710);
   U18050 : AOI221_X1 port map( B1 => n23276, B2 => n20937, C1 => n22494, C2 =>
                           n21677, A => n24710, ZN => n24711);
   U18051 : NAND4_X1 port map( A1 => n24712, A2 => n24713, A3 => n24711, A4 => 
                           n24714, ZN => n3296);
   U18052 : NAND2_X1 port map( A1 => n17907, A2 => n17908, ZN => n24716);
   U18053 : AOI21_X1 port map( B1 => n17911, B2 => n17912, A => n23197, ZN => 
                           n24715);
   U18054 : AOI221_X1 port map( B1 => n23213, B2 => n21901, C1 => n23205, C2 =>
                           n24716, A => n24715, ZN => n24720);
   U18055 : AOI222_X1 port map( A1 => n23237, A2 => n21344, B1 => n23229, B2 =>
                           n21020, C1 => n23221, C2 => n20827, ZN => n24719);
   U18056 : OAI222_X1 port map( A1 => n20455, A2 => n23261, B1 => n20583, B2 =>
                           n23253, C1 => n20519, C2 => n23245, ZN => n24717);
   U18057 : NOR4_X1 port map( A1 => n24717, A2 => n17916, A3 => n17903, A4 => 
                           n17904, ZN => n24718);
   U18058 : AND3_X1 port map( A1 => n24720, A2 => n24719, A3 => n24718, ZN => 
                           n24721);
   U18059 : OAI22_X1 port map( A1 => n19175, A2 => n22976, B1 => n19303, B2 => 
                           n22650, ZN => n24723);
   U18060 : AOI221_X1 port map( B1 => n22911, B2 => n22086, C1 => n22804, C2 =>
                           n21209, A => n24723, ZN => n24729);
   U18061 : OAI222_X1 port map( A1 => n18983, A2 => n22954, B1 => n19239, B2 =>
                           n22967, C1 => n19111, C2 => n22639, ZN => n24724);
   U18062 : AOI221_X1 port map( B1 => n22801, B2 => n22042, C1 => n22960, C2 =>
                           n21274, A => n24724, ZN => n24728);
   U18063 : OAI22_X1 port map( A1 => n23270, A2 => n24725, B1 => n18727, B2 => 
                           n22947, ZN => n24726);
   U18064 : AOI221_X1 port map( B1 => n23276, B2 => n20956, C1 => n22494, C2 =>
                           n21764, A => n24726, ZN => n24727);
   U18065 : NAND4_X1 port map( A1 => n24727, A2 => n24730, A3 => n24728, A4 => 
                           n24729, ZN => n3297);
   U18066 : NAND2_X1 port map( A1 => n17880, A2 => n17881, ZN => n24732);
   U18067 : AOI21_X1 port map( B1 => n17884, B2 => n17885, A => n23197, ZN => 
                           n24731);
   U18068 : AOI221_X1 port map( B1 => n23213, B2 => n21869, C1 => n23205, C2 =>
                           n24732, A => n24731, ZN => n24736);
   U18069 : AOI222_X1 port map( A1 => n23237, A2 => n21312, B1 => n23229, B2 =>
                           n20988, C1 => n23221, C2 => n20795, ZN => n24735);
   U18070 : OAI222_X1 port map( A1 => n20432, A2 => n23261, B1 => n20560, B2 =>
                           n23253, C1 => n20496, C2 => n23245, ZN => n24733);
   U18071 : NOR4_X1 port map( A1 => n24733, A2 => n17889, A3 => n17876, A4 => 
                           n17877, ZN => n24734);
   U18072 : AND3_X1 port map( A1 => n24736, A2 => n24735, A3 => n24734, ZN => 
                           n24737);
   U18073 : OAI222_X1 port map( A1 => n19536, A2 => n22652, B1 => n24737, B2 =>
                           n22800, C1 => n19664, C2 => n22518, ZN => n24738);
   U18074 : AOI221_X1 port map( B1 => n22923, B2 => n22106, C1 => n22969, C2 =>
                           n21119, A => n24738, ZN => n24746);
   U18075 : OAI22_X1 port map( A1 => n19152, A2 => n22980, B1 => n19280, B2 => 
                           n22646, ZN => n24739);
   U18076 : AOI221_X1 port map( B1 => n22915, B2 => n22067, C1 => n22805, C2 =>
                           n21161, A => n24739, ZN => n24745);
   U18077 : OAI222_X1 port map( A1 => n18960, A2 => n22955, B1 => n19216, B2 =>
                           n22964, C1 => n19088, C2 => n22639, ZN => n24740);
   U18078 : AOI221_X1 port map( B1 => n25391, B2 => n22159, C1 => n22959, C2 =>
                           n21235, A => n24740, ZN => n24744);
   U18079 : OAI22_X1 port map( A1 => n23269, A2 => n24741, B1 => n18704, B2 => 
                           n22943, ZN => n24742);
   U18080 : AOI221_X1 port map( B1 => n23276, B2 => n20924, C1 => n22494, C2 =>
                           n21664, A => n24742, ZN => n24743);
   U18081 : NAND4_X1 port map( A1 => n24744, A2 => n24745, A3 => n24743, A4 => 
                           n24746, ZN => n3298);
   U18082 : NAND2_X1 port map( A1 => n17853, A2 => n17854, ZN => n24748);
   U18083 : AOI21_X1 port map( B1 => n17857, B2 => n17858, A => n23198, ZN => 
                           n24747);
   U18084 : AOI221_X1 port map( B1 => n23214, B2 => n21847, C1 => n23206, C2 =>
                           n24748, A => n24747, ZN => n24752);
   U18085 : AOI222_X1 port map( A1 => n23238, A2 => n21290, B1 => n23230, B2 =>
                           n20966, C1 => n23222, C2 => n20773, ZN => n24751);
   U18086 : OAI222_X1 port map( A1 => n20456, A2 => n23262, B1 => n20584, B2 =>
                           n23254, C1 => n20520, C2 => n23246, ZN => n24749);
   U18087 : NOR4_X1 port map( A1 => n24749, A2 => n17862, A3 => n17849, A4 => 
                           n17850, ZN => n24750);
   U18088 : AND3_X1 port map( A1 => n24752, A2 => n24751, A3 => n24750, ZN => 
                           n24753);
   U18089 : OAI222_X1 port map( A1 => n19560, A2 => n22652, B1 => n24753, B2 =>
                           n22798, C1 => n19688, C2 => n22518, ZN => n24754);
   U18090 : AOI221_X1 port map( B1 => n22921, B2 => n22107, C1 => n22975, C2 =>
                           n21097, A => n24754, ZN => n24762);
   U18091 : OAI22_X1 port map( A1 => n19176, A2 => n22979, B1 => n19304, B2 => 
                           n22633, ZN => n24755);
   U18092 : OAI222_X1 port map( A1 => n18984, A2 => n22953, B1 => n19240, B2 =>
                           n22964, C1 => n19112, C2 => n22637, ZN => n24756);
   U18093 : AOI221_X1 port map( B1 => n25391, B2 => n22160, C1 => n22958, C2 =>
                           n21213, A => n24756, ZN => n24760);
   U18094 : OAI22_X1 port map( A1 => n25394, A2 => n24757, B1 => n18728, B2 => 
                           n22947, ZN => n24758);
   U18095 : NAND4_X1 port map( A1 => n24760, A2 => n24761, A3 => n24759, A4 => 
                           n24762, ZN => n3299);
   U18096 : NAND2_X1 port map( A1 => n17826, A2 => n17827, ZN => n24764);
   U18097 : AOI21_X1 port map( B1 => n17830, B2 => n17831, A => n23198, ZN => 
                           n24763);
   U18098 : AOI221_X1 port map( B1 => n23214, B2 => n21883, C1 => n23206, C2 =>
                           n24764, A => n24763, ZN => n24768);
   U18099 : AOI222_X1 port map( A1 => n23238, A2 => n21326, B1 => n23230, B2 =>
                           n21002, C1 => n23222, C2 => n20809, ZN => n24767);
   U18100 : OAI222_X1 port map( A1 => n20431, A2 => n23262, B1 => n20559, B2 =>
                           n23254, C1 => n20495, C2 => n23246, ZN => n24765);
   U18101 : NOR4_X1 port map( A1 => n24765, A2 => n17835, A3 => n17822, A4 => 
                           n17823, ZN => n24766);
   U18102 : AND3_X1 port map( A1 => n24768, A2 => n24767, A3 => n24766, ZN => 
                           n24769);
   U18103 : OAI222_X1 port map( A1 => n19535, A2 => n22652, B1 => n24769, B2 =>
                           n22799, C1 => n19663, C2 => n22517, ZN => n24770);
   U18104 : AOI221_X1 port map( B1 => n22523, B2 => n22108, C1 => n22975, C2 =>
                           n21132, A => n24770, ZN => n24778);
   U18105 : OAI22_X1 port map( A1 => n19151, A2 => n22978, B1 => n19279, B2 => 
                           n22645, ZN => n24771);
   U18106 : OAI222_X1 port map( A1 => n18959, A2 => n22953, B1 => n19215, B2 =>
                           n22967, C1 => n19087, C2 => n22636, ZN => n24772);
   U18107 : AOI221_X1 port map( B1 => n22801, B2 => n22043, C1 => n22958, C2 =>
                           n21250, A => n24772, ZN => n24776);
   U18108 : OAI22_X1 port map( A1 => n25394, A2 => n24773, B1 => n18703, B2 => 
                           n22943, ZN => n24774);
   U18109 : AOI221_X1 port map( B1 => n23277, B2 => n20938, C1 => n22494, C2 =>
                           n21678, A => n24774, ZN => n24775);
   U18110 : NAND4_X1 port map( A1 => n24775, A2 => n24777, A3 => n24776, A4 => 
                           n24778, ZN => n3300);
   U18111 : NAND2_X1 port map( A1 => n17799, A2 => n17800, ZN => n24780);
   U18112 : AOI21_X1 port map( B1 => n17803, B2 => n17804, A => n23198, ZN => 
                           n24779);
   U18113 : AOI221_X1 port map( B1 => n23214, B2 => n21848, C1 => n23206, C2 =>
                           n24780, A => n24779, ZN => n24784);
   U18114 : AOI222_X1 port map( A1 => n23238, A2 => n21291, B1 => n23230, B2 =>
                           n20967, C1 => n23222, C2 => n20774, ZN => n24783);
   U18115 : OAI222_X1 port map( A1 => n20457, A2 => n23262, B1 => n20585, B2 =>
                           n23254, C1 => n20521, C2 => n23246, ZN => n24781);
   U18116 : NOR4_X1 port map( A1 => n24781, A2 => n17808, A3 => n17795, A4 => 
                           n17796, ZN => n24782);
   U18117 : AND3_X1 port map( A1 => n24784, A2 => n24783, A3 => n24782, ZN => 
                           n24785);
   U18118 : OAI222_X1 port map( A1 => n19561, A2 => n22652, B1 => n24785, B2 =>
                           n22798, C1 => n19689, C2 => n22518, ZN => n24786);
   U18119 : AOI221_X1 port map( B1 => n22522, B2 => n22109, C1 => n22974, C2 =>
                           n21098, A => n24786, ZN => n24794);
   U18120 : OAI22_X1 port map( A1 => n19177, A2 => n22979, B1 => n19305, B2 => 
                           n22641, ZN => n24787);
   U18121 : OAI222_X1 port map( A1 => n18985, A2 => n22951, B1 => n19241, B2 =>
                           n22964, C1 => n19113, C2 => n22636, ZN => n24788);
   U18122 : AOI221_X1 port map( B1 => n22801, B2 => n22044, C1 => n22959, C2 =>
                           n21214, A => n24788, ZN => n24792);
   U18123 : OAI22_X1 port map( A1 => n23270, A2 => n24789, B1 => n18729, B2 => 
                           n22944, ZN => n24790);
   U18124 : AOI221_X1 port map( B1 => n23277, B2 => n20903, C1 => n22494, C2 =>
                           n21643, A => n24790, ZN => n24791);
   U18125 : NAND4_X1 port map( A1 => n24791, A2 => n24793, A3 => n24792, A4 => 
                           n24794, ZN => n3301);
   U18126 : NAND2_X1 port map( A1 => n17772, A2 => n17773, ZN => n24796);
   U18127 : AOI21_X1 port map( B1 => n17776, B2 => n17777, A => n23198, ZN => 
                           n24795);
   U18128 : AOI221_X1 port map( B1 => n23214, B2 => n21870, C1 => n23206, C2 =>
                           n24796, A => n24795, ZN => n24800);
   U18129 : AOI222_X1 port map( A1 => n23238, A2 => n21313, B1 => n23230, B2 =>
                           n20989, C1 => n23222, C2 => n20796, ZN => n24799);
   U18130 : OAI222_X1 port map( A1 => n20430, A2 => n23262, B1 => n20558, B2 =>
                           n23254, C1 => n20494, C2 => n23246, ZN => n24797);
   U18131 : NOR4_X1 port map( A1 => n24797, A2 => n17781, A3 => n17768, A4 => 
                           n17769, ZN => n24798);
   U18132 : AND3_X1 port map( A1 => n24800, A2 => n24799, A3 => n24798, ZN => 
                           n24801);
   U18133 : OAI222_X1 port map( A1 => n19534, A2 => n22935, B1 => n24801, B2 =>
                           n22800, C1 => n19662, C2 => n22520, ZN => n24802);
   U18134 : AOI221_X1 port map( B1 => n22921, B2 => n22110, C1 => n22975, C2 =>
                           n21120, A => n24802, ZN => n24810);
   U18135 : OAI22_X1 port map( A1 => n19150, A2 => n22978, B1 => n19278, B2 => 
                           n22630, ZN => n24803);
   U18136 : AOI221_X1 port map( B1 => n22916, B2 => n22068, C1 => n22812, C2 =>
                           n21162, A => n24803, ZN => n24809);
   U18137 : OAI222_X1 port map( A1 => n18958, A2 => n22955, B1 => n19214, B2 =>
                           n22965, C1 => n19086, C2 => n22636, ZN => n24804);
   U18138 : AOI221_X1 port map( B1 => n22801, B2 => n22045, C1 => n22960, C2 =>
                           n21236, A => n24804, ZN => n24808);
   U18139 : OAI22_X1 port map( A1 => n23269, A2 => n24805, B1 => n18702, B2 => 
                           n22943, ZN => n24806);
   U18140 : AOI221_X1 port map( B1 => n23277, B2 => n20925, C1 => n22494, C2 =>
                           n21665, A => n24806, ZN => n24807);
   U18141 : NAND4_X1 port map( A1 => n24807, A2 => n24809, A3 => n24808, A4 => 
                           n24810, ZN => n3302);
   U18142 : NAND2_X1 port map( A1 => n17745, A2 => n17746, ZN => n24812);
   U18143 : AOI21_X1 port map( B1 => n17749, B2 => n17750, A => n23198, ZN => 
                           n24811);
   U18144 : AOI221_X1 port map( B1 => n23214, B2 => n21884, C1 => n23206, C2 =>
                           n24812, A => n24811, ZN => n24816);
   U18145 : AOI222_X1 port map( A1 => n23238, A2 => n21327, B1 => n23230, B2 =>
                           n21003, C1 => n23222, C2 => n20810, ZN => n24815);
   U18146 : OAI222_X1 port map( A1 => n20458, A2 => n23262, B1 => n20586, B2 =>
                           n23254, C1 => n20522, C2 => n23246, ZN => n24813);
   U18147 : NOR4_X1 port map( A1 => n24813, A2 => n17754, A3 => n17741, A4 => 
                           n17742, ZN => n24814);
   U18148 : AND3_X1 port map( A1 => n24816, A2 => n24815, A3 => n24814, ZN => 
                           n24817);
   U18149 : OAI222_X1 port map( A1 => n19562, A2 => n22937, B1 => n24817, B2 =>
                           n22799, C1 => n19690, C2 => n22517, ZN => n24818);
   U18150 : AOI221_X1 port map( B1 => n22522, B2 => n22111, C1 => n22975, C2 =>
                           n21133, A => n24818, ZN => n24826);
   U18151 : OAI22_X1 port map( A1 => n19178, A2 => n22977, B1 => n19306, B2 => 
                           n22644, ZN => n24819);
   U18152 : OAI222_X1 port map( A1 => n18986, A2 => n22954, B1 => n19242, B2 =>
                           n22967, C1 => n19114, C2 => n22637, ZN => n24820);
   U18153 : AOI221_X1 port map( B1 => n22801, B2 => n22046, C1 => n22959, C2 =>
                           n21251, A => n24820, ZN => n24824);
   U18154 : OAI22_X1 port map( A1 => n23269, A2 => n24821, B1 => n18730, B2 => 
                           n22944, ZN => n24822);
   U18155 : AOI221_X1 port map( B1 => n23277, B2 => n20939, C1 => n22494, C2 =>
                           n21679, A => n24822, ZN => n24823);
   U18156 : NAND4_X1 port map( A1 => n24823, A2 => n24825, A3 => n24824, A4 => 
                           n24826, ZN => n3303);
   U18157 : NAND2_X1 port map( A1 => n17718, A2 => n17719, ZN => n24828);
   U18158 : AOI21_X1 port map( B1 => n17722, B2 => n17723, A => n23198, ZN => 
                           n24827);
   U18159 : AOI221_X1 port map( B1 => n23214, B2 => n21871, C1 => n23206, C2 =>
                           n24828, A => n24827, ZN => n24832);
   U18160 : AOI222_X1 port map( A1 => n23238, A2 => n21314, B1 => n23230, B2 =>
                           n20990, C1 => n23222, C2 => n20797, ZN => n24831);
   U18161 : OAI222_X1 port map( A1 => n20429, A2 => n23262, B1 => n20557, B2 =>
                           n23254, C1 => n20493, C2 => n23246, ZN => n24829);
   U18162 : NOR4_X1 port map( A1 => n24829, A2 => n17727, A3 => n17714, A4 => 
                           n17715, ZN => n24830);
   U18163 : AND3_X1 port map( A1 => n24832, A2 => n24831, A3 => n24830, ZN => 
                           n24833);
   U18164 : OAI222_X1 port map( A1 => n19533, A2 => n22652, B1 => n24833, B2 =>
                           n22800, C1 => n19661, C2 => n22519, ZN => n24834);
   U18165 : AOI221_X1 port map( B1 => n22922, B2 => n22112, C1 => n22975, C2 =>
                           n21121, A => n24834, ZN => n24842);
   U18166 : OAI22_X1 port map( A1 => n19149, A2 => n22976, B1 => n19277, B2 => 
                           n22647, ZN => n24835);
   U18167 : OAI222_X1 port map( A1 => n18957, A2 => n22953, B1 => n19213, B2 =>
                           n22966, C1 => n19085, C2 => n22638, ZN => n24836);
   U18168 : AOI221_X1 port map( B1 => n22801, B2 => n22047, C1 => n22957, C2 =>
                           n21237, A => n24836, ZN => n24840);
   U18169 : OAI22_X1 port map( A1 => n25394, A2 => n24837, B1 => n18701, B2 => 
                           n22945, ZN => n24838);
   U18170 : AOI221_X1 port map( B1 => n23277, B2 => n20926, C1 => n22494, C2 =>
                           n21666, A => n24838, ZN => n24839);
   U18171 : NAND4_X1 port map( A1 => n24839, A2 => n24841, A3 => n24840, A4 => 
                           n24842, ZN => n3304);
   U18172 : NAND2_X1 port map( A1 => n17691, A2 => n17692, ZN => n24844);
   U18173 : AOI21_X1 port map( B1 => n17695, B2 => n17696, A => n23198, ZN => 
                           n24843);
   U18174 : AOI221_X1 port map( B1 => n23214, B2 => n21872, C1 => n23206, C2 =>
                           n24844, A => n24843, ZN => n24848);
   U18175 : AOI222_X1 port map( A1 => n23238, A2 => n21315, B1 => n23230, B2 =>
                           n20991, C1 => n23222, C2 => n20798, ZN => n24847);
   U18176 : OAI222_X1 port map( A1 => n20459, A2 => n23262, B1 => n20587, B2 =>
                           n23254, C1 => n20523, C2 => n23246, ZN => n24845);
   U18177 : NOR4_X1 port map( A1 => n24845, A2 => n17700, A3 => n17687, A4 => 
                           n17688, ZN => n24846);
   U18178 : AND3_X1 port map( A1 => n24848, A2 => n24847, A3 => n24846, ZN => 
                           n24849);
   U18179 : OAI222_X1 port map( A1 => n19563, A2 => n22934, B1 => n24849, B2 =>
                           n22800, C1 => n19691, C2 => n22516, ZN => n24850);
   U18180 : AOI221_X1 port map( B1 => n22923, B2 => n22113, C1 => n22975, C2 =>
                           n21122, A => n24850, ZN => n24858);
   U18181 : OAI22_X1 port map( A1 => n19179, A2 => n22977, B1 => n19307, B2 => 
                           n22642, ZN => n24851);
   U18182 : OAI222_X1 port map( A1 => n18987, A2 => n22952, B1 => n19243, B2 =>
                           n22967, C1 => n19115, C2 => n22637, ZN => n24852);
   U18183 : AOI221_X1 port map( B1 => n22801, B2 => n22048, C1 => n22958, C2 =>
                           n21238, A => n24852, ZN => n24856);
   U18184 : OAI22_X1 port map( A1 => n23270, A2 => n24853, B1 => n18731, B2 => 
                           n22946, ZN => n24854);
   U18185 : AOI221_X1 port map( B1 => n23277, B2 => n20927, C1 => n22494, C2 =>
                           n21667, A => n24854, ZN => n24855);
   U18186 : NAND4_X1 port map( A1 => n24855, A2 => n24857, A3 => n24856, A4 => 
                           n24858, ZN => n3305);
   U18187 : NAND2_X1 port map( A1 => n17664, A2 => n17665, ZN => n24860);
   U18188 : AOI21_X1 port map( B1 => n17668, B2 => n17669, A => n23198, ZN => 
                           n24859);
   U18189 : AOI221_X1 port map( B1 => n23214, B2 => n21873, C1 => n23206, C2 =>
                           n24860, A => n24859, ZN => n24864);
   U18190 : AOI222_X1 port map( A1 => n23238, A2 => n21316, B1 => n23230, B2 =>
                           n20992, C1 => n23222, C2 => n20799, ZN => n24863);
   U18191 : OAI222_X1 port map( A1 => n20428, A2 => n23262, B1 => n20556, B2 =>
                           n23254, C1 => n20492, C2 => n23246, ZN => n24861);
   U18192 : NOR4_X1 port map( A1 => n24861, A2 => n17673, A3 => n17660, A4 => 
                           n17661, ZN => n24862);
   U18193 : AND3_X1 port map( A1 => n24864, A2 => n24863, A3 => n24862, ZN => 
                           n24865);
   U18194 : OAI222_X1 port map( A1 => n19532, A2 => n22935, B1 => n24865, B2 =>
                           n22800, C1 => n19660, C2 => n22518, ZN => n24866);
   U18195 : AOI221_X1 port map( B1 => n22523, B2 => n22114, C1 => n22975, C2 =>
                           n21123, A => n24866, ZN => n24874);
   U18196 : OAI22_X1 port map( A1 => n19148, A2 => n22978, B1 => n19276, B2 => 
                           n22634, ZN => n24867);
   U18197 : AOI221_X1 port map( B1 => n22919, B2 => n22069, C1 => n22809, C2 =>
                           n21163, A => n24867, ZN => n24873);
   U18198 : OAI222_X1 port map( A1 => n18956, A2 => n22952, B1 => n19212, B2 =>
                           n22965, C1 => n19084, C2 => n22637, ZN => n24868);
   U18199 : AOI221_X1 port map( B1 => n22801, B2 => n22049, C1 => n22959, C2 =>
                           n21239, A => n24868, ZN => n24872);
   U18200 : OAI22_X1 port map( A1 => n23269, A2 => n24869, B1 => n18700, B2 => 
                           n22947, ZN => n24870);
   U18201 : AOI221_X1 port map( B1 => n23277, B2 => n20928, C1 => n22494, C2 =>
                           n21668, A => n24870, ZN => n24871);
   U18202 : NAND4_X1 port map( A1 => n24871, A2 => n24873, A3 => n24872, A4 => 
                           n24874, ZN => n3306);
   U18203 : NAND2_X1 port map( A1 => n17637, A2 => n17638, ZN => n24876);
   U18204 : AOI21_X1 port map( B1 => n17641, B2 => n17642, A => n23198, ZN => 
                           n24875);
   U18205 : AOI221_X1 port map( B1 => n23214, B2 => n21904, C1 => n23206, C2 =>
                           n24876, A => n24875, ZN => n24880);
   U18206 : AOI222_X1 port map( A1 => n23238, A2 => n21347, B1 => n23230, B2 =>
                           n21023, C1 => n23222, C2 => n20830, ZN => n24879);
   U18207 : OAI222_X1 port map( A1 => n20460, A2 => n23262, B1 => n20588, B2 =>
                           n23254, C1 => n20524, C2 => n23246, ZN => n24877);
   U18208 : NOR4_X1 port map( A1 => n24877, A2 => n17646, A3 => n17633, A4 => 
                           n17634, ZN => n24878);
   U18209 : AND3_X1 port map( A1 => n24880, A2 => n24879, A3 => n24878, ZN => 
                           n24881);
   U18210 : OAI222_X1 port map( A1 => n19564, A2 => n22934, B1 => n24881, B2 =>
                           n22799, C1 => n19692, C2 => n22519, ZN => n24882);
   U18211 : OAI22_X1 port map( A1 => n19180, A2 => n22980, B1 => n19308, B2 => 
                           n22649, ZN => n24883);
   U18212 : AOI221_X1 port map( B1 => n22914, B2 => n22070, C1 => n22806, C2 =>
                           n21275, A => n24883, ZN => n24889);
   U18213 : OAI222_X1 port map( A1 => n18988, A2 => n22955, B1 => n19244, B2 =>
                           n22966, C1 => n19116, C2 => n22639, ZN => n24884);
   U18214 : AOI221_X1 port map( B1 => n22801, B2 => n22050, C1 => n22960, C2 =>
                           n21281, A => n24884, ZN => n24888);
   U18215 : OAI22_X1 port map( A1 => n25394, A2 => n24885, B1 => n18732, B2 => 
                           n22944, ZN => n24886);
   U18216 : AOI221_X1 port map( B1 => n23277, B2 => n20959, C1 => n22494, C2 =>
                           n21832, A => n24886, ZN => n24887);
   U18217 : NAND4_X1 port map( A1 => n24887, A2 => n24889, A3 => n24888, A4 => 
                           n24890, ZN => n3307);
   U18218 : NAND2_X1 port map( A1 => n17610, A2 => n17611, ZN => n24892);
   U18219 : AOI21_X1 port map( B1 => n17614, B2 => n17615, A => n23198, ZN => 
                           n24891);
   U18220 : AOI221_X1 port map( B1 => n23214, B2 => n21849, C1 => n23206, C2 =>
                           n24892, A => n24891, ZN => n24896);
   U18221 : AOI222_X1 port map( A1 => n23238, A2 => n21292, B1 => n23230, B2 =>
                           n20968, C1 => n23222, C2 => n20775, ZN => n24895);
   U18222 : OAI222_X1 port map( A1 => n20427, A2 => n23262, B1 => n20555, B2 =>
                           n23254, C1 => n20491, C2 => n23246, ZN => n24893);
   U18223 : NOR4_X1 port map( A1 => n24893, A2 => n17619, A3 => n17606, A4 => 
                           n17607, ZN => n24894);
   U18224 : AND3_X1 port map( A1 => n24896, A2 => n24895, A3 => n24894, ZN => 
                           n24897);
   U18225 : OAI222_X1 port map( A1 => n19531, A2 => n22934, B1 => n24897, B2 =>
                           n22798, C1 => n19659, C2 => n22521, ZN => n24898);
   U18226 : AOI221_X1 port map( B1 => n22522, B2 => n22115, C1 => n22975, C2 =>
                           n21099, A => n24898, ZN => n24906);
   U18227 : OAI22_X1 port map( A1 => n19147, A2 => n22979, B1 => n19275, B2 => 
                           n22646, ZN => n24899);
   U18228 : AOI221_X1 port map( B1 => n22916, B2 => n22071, C1 => n22810, C2 =>
                           n21153, A => n24899, ZN => n24905);
   U18229 : OAI222_X1 port map( A1 => n18955, A2 => n22952, B1 => n19211, B2 =>
                           n22966, C1 => n19083, C2 => n22637, ZN => n24900);
   U18230 : AOI221_X1 port map( B1 => n22801, B2 => n22051, C1 => n22961, C2 =>
                           n21215, A => n24900, ZN => n24904);
   U18231 : OAI22_X1 port map( A1 => n23270, A2 => n24901, B1 => n18699, B2 => 
                           n22945, ZN => n24902);
   U18232 : AOI221_X1 port map( B1 => n23277, B2 => n20904, C1 => n22494, C2 =>
                           n21644, A => n24902, ZN => n24903);
   U18233 : NAND4_X1 port map( A1 => n24903, A2 => n24905, A3 => n24904, A4 => 
                           n24906, ZN => n3308);
   U18234 : NAND2_X1 port map( A1 => n17583, A2 => n17584, ZN => n24908);
   U18235 : AOI21_X1 port map( B1 => n17587, B2 => n17588, A => n23198, ZN => 
                           n24907);
   U18236 : AOI221_X1 port map( B1 => n23214, B2 => n21885, C1 => n23206, C2 =>
                           n24908, A => n24907, ZN => n24912);
   U18237 : AOI222_X1 port map( A1 => n23238, A2 => n21328, B1 => n23230, B2 =>
                           n21004, C1 => n23222, C2 => n20811, ZN => n24911);
   U18238 : OAI222_X1 port map( A1 => n20461, A2 => n23262, B1 => n20589, B2 =>
                           n23254, C1 => n20525, C2 => n23246, ZN => n24909);
   U18239 : NOR4_X1 port map( A1 => n24909, A2 => n17592, A3 => n17579, A4 => 
                           n17580, ZN => n24910);
   U18240 : AND3_X1 port map( A1 => n24912, A2 => n24911, A3 => n24910, ZN => 
                           n24913);
   U18241 : OAI222_X1 port map( A1 => n19565, A2 => n22934, B1 => n24913, B2 =>
                           n22799, C1 => n19693, C2 => n22520, ZN => n24914);
   U18242 : AOI221_X1 port map( B1 => n22922, B2 => n22116, C1 => n22975, C2 =>
                           n21134, A => n24914, ZN => n24922);
   U18243 : OAI22_X1 port map( A1 => n19181, A2 => n22978, B1 => n19309, B2 => 
                           n22630, ZN => n24915);
   U18244 : AOI221_X1 port map( B1 => n22920, B2 => n22072, C1 => n22804, C2 =>
                           n21168, A => n24915, ZN => n24921);
   U18245 : OAI222_X1 port map( A1 => n18989, A2 => n22951, B1 => n19245, B2 =>
                           n22964, C1 => n19117, C2 => n22638, ZN => n24916);
   U18246 : AOI221_X1 port map( B1 => n25391, B2 => n22161, C1 => n22957, C2 =>
                           n21252, A => n24916, ZN => n24920);
   U18247 : OAI22_X1 port map( A1 => n23269, A2 => n24917, B1 => n18733, B2 => 
                           n22943, ZN => n24918);
   U18248 : AOI221_X1 port map( B1 => n23277, B2 => n20940, C1 => n22494, C2 =>
                           n21680, A => n24918, ZN => n24919);
   U18249 : NAND4_X1 port map( A1 => n24920, A2 => n24921, A3 => n24919, A4 => 
                           n24922, ZN => n3309);
   U18250 : NAND2_X1 port map( A1 => n17556, A2 => n17557, ZN => n24924);
   U18251 : AOI21_X1 port map( B1 => n17560, B2 => n17561, A => n23198, ZN => 
                           n24923);
   U18252 : AOI221_X1 port map( B1 => n23214, B2 => n21850, C1 => n23206, C2 =>
                           n24924, A => n24923, ZN => n24928);
   U18253 : AOI222_X1 port map( A1 => n23238, A2 => n21293, B1 => n23230, B2 =>
                           n20969, C1 => n23222, C2 => n20776, ZN => n24927);
   U18254 : OAI222_X1 port map( A1 => n20426, A2 => n23262, B1 => n20554, B2 =>
                           n23254, C1 => n20490, C2 => n23246, ZN => n24925);
   U18255 : NOR4_X1 port map( A1 => n24925, A2 => n17565, A3 => n17552, A4 => 
                           n17553, ZN => n24926);
   U18256 : AND3_X1 port map( A1 => n24928, A2 => n24927, A3 => n24926, ZN => 
                           n24929);
   U18257 : OAI222_X1 port map( A1 => n19530, A2 => n22936, B1 => n24929, B2 =>
                           n22798, C1 => n19658, C2 => n22517, ZN => n24930);
   U18258 : AOI221_X1 port map( B1 => n22922, B2 => n22117, C1 => n22971, C2 =>
                           n21100, A => n24930, ZN => n24938);
   U18259 : OAI22_X1 port map( A1 => n19146, A2 => n22976, B1 => n19274, B2 => 
                           n22646, ZN => n24931);
   U18260 : AOI221_X1 port map( B1 => n22920, B2 => n22073, C1 => n22805, C2 =>
                           n21154, A => n24931, ZN => n24937);
   U18261 : OAI222_X1 port map( A1 => n18954, A2 => n22951, B1 => n19210, B2 =>
                           n22967, C1 => n19082, C2 => n22636, ZN => n24932);
   U18262 : AOI221_X1 port map( B1 => n25391, B2 => n22162, C1 => n22961, C2 =>
                           n21216, A => n24932, ZN => n24936);
   U18263 : OAI22_X1 port map( A1 => n25394, A2 => n24933, B1 => n18698, B2 => 
                           n22944, ZN => n24934);
   U18264 : AOI221_X1 port map( B1 => n23277, B2 => n20905, C1 => n22494, C2 =>
                           n21645, A => n24934, ZN => n24935);
   U18265 : NAND4_X1 port map( A1 => n24936, A2 => n24937, A3 => n24935, A4 => 
                           n24938, ZN => n3310);
   U18266 : NAND2_X1 port map( A1 => n17529, A2 => n17530, ZN => n24940);
   U18267 : AOI21_X1 port map( B1 => n17533, B2 => n17534, A => n23199, ZN => 
                           n24939);
   U18268 : AOI221_X1 port map( B1 => n23215, B2 => n21905, C1 => n23207, C2 =>
                           n24940, A => n24939, ZN => n24944);
   U18269 : AOI222_X1 port map( A1 => n23239, A2 => n21348, B1 => n23231, B2 =>
                           n21024, C1 => n23223, C2 => n20831, ZN => n24943);
   U18270 : OAI222_X1 port map( A1 => n20462, A2 => n23263, B1 => n20590, B2 =>
                           n23255, C1 => n20526, C2 => n23247, ZN => n24941);
   U18271 : NOR4_X1 port map( A1 => n24941, A2 => n17538, A3 => n17525, A4 => 
                           n17526, ZN => n24942);
   U18272 : AND3_X1 port map( A1 => n24944, A2 => n24943, A3 => n24942, ZN => 
                           n24945);
   U18273 : OAI222_X1 port map( A1 => n19566, A2 => n22936, B1 => n24945, B2 =>
                           n22799, C1 => n19694, C2 => n22518, ZN => n24946);
   U18274 : OAI22_X1 port map( A1 => n19182, A2 => n22977, B1 => n19310, B2 => 
                           n22631, ZN => n24947);
   U18275 : AOI221_X1 port map( B1 => n22920, B2 => n22074, C1 => n22809, C2 =>
                           n21276, A => n24947, ZN => n24953);
   U18276 : OAI222_X1 port map( A1 => n18990, A2 => n22951, B1 => n19246, B2 =>
                           n22964, C1 => n19118, C2 => n22636, ZN => n24948);
   U18277 : AOI221_X1 port map( B1 => n25391, B2 => n22163, C1 => n22962, C2 =>
                           n21282, A => n24948, ZN => n24952);
   U18278 : OAI22_X1 port map( A1 => n25394, A2 => n24949, B1 => n18734, B2 => 
                           n22945, ZN => n24950);
   U18279 : AOI221_X1 port map( B1 => n23278, B2 => n20960, C1 => n22494, C2 =>
                           n21833, A => n24950, ZN => n24951);
   U18280 : NAND4_X1 port map( A1 => n24952, A2 => n24953, A3 => n24951, A4 => 
                           n24954, ZN => n3311);
   U18281 : NAND2_X1 port map( A1 => n17502, A2 => n17503, ZN => n24956);
   U18282 : AOI21_X1 port map( B1 => n17506, B2 => n17507, A => n23199, ZN => 
                           n24955);
   U18283 : AOI221_X1 port map( B1 => n23215, B2 => n21906, C1 => n23207, C2 =>
                           n24956, A => n24955, ZN => n24960);
   U18284 : AOI222_X1 port map( A1 => n23239, A2 => n21349, B1 => n23231, B2 =>
                           n21025, C1 => n23223, C2 => n20832, ZN => n24959);
   U18285 : OAI222_X1 port map( A1 => n20425, A2 => n23263, B1 => n20553, B2 =>
                           n23255, C1 => n20489, C2 => n23247, ZN => n24957);
   U18286 : NOR4_X1 port map( A1 => n24957, A2 => n17511, A3 => n17498, A4 => 
                           n17499, ZN => n24958);
   U18287 : AND3_X1 port map( A1 => n24960, A2 => n24959, A3 => n24958, ZN => 
                           n24961);
   U18288 : OAI222_X1 port map( A1 => n19529, A2 => n22937, B1 => n24961, B2 =>
                           n22799, C1 => n19657, C2 => n22517, ZN => n24962);
   U18289 : OAI22_X1 port map( A1 => n19145, A2 => n22977, B1 => n19273, B2 => 
                           n22647, ZN => n24963);
   U18290 : AOI221_X1 port map( B1 => n22920, B2 => n22075, C1 => n22804, C2 =>
                           n21277, A => n24963, ZN => n24969);
   U18291 : OAI222_X1 port map( A1 => n18953, A2 => n22955, B1 => n19209, B2 =>
                           n22968, C1 => n19081, C2 => n22635, ZN => n24964);
   U18292 : AOI221_X1 port map( B1 => n25391, B2 => n22164, C1 => n22962, C2 =>
                           n21283, A => n24964, ZN => n24968);
   U18293 : OAI22_X1 port map( A1 => n23269, A2 => n24965, B1 => n18697, B2 => 
                           n22945, ZN => n24966);
   U18294 : AOI221_X1 port map( B1 => n23278, B2 => n20961, C1 => n22494, C2 =>
                           n21834, A => n24966, ZN => n24967);
   U18295 : NAND4_X1 port map( A1 => n24968, A2 => n24969, A3 => n24967, A4 => 
                           n24970, ZN => n3312);
   U18296 : NAND2_X1 port map( A1 => n17475, A2 => n17476, ZN => n24972);
   U18297 : AOI21_X1 port map( B1 => n17479, B2 => n17480, A => n23199, ZN => 
                           n24971);
   U18298 : AOI221_X1 port map( B1 => n23215, B2 => n21874, C1 => n23207, C2 =>
                           n24972, A => n24971, ZN => n24976);
   U18299 : AOI222_X1 port map( A1 => n23239, A2 => n21317, B1 => n23231, B2 =>
                           n20993, C1 => n23223, C2 => n20800, ZN => n24975);
   U18300 : OAI222_X1 port map( A1 => n20463, A2 => n23263, B1 => n20591, B2 =>
                           n23255, C1 => n20527, C2 => n23247, ZN => n24973);
   U18301 : NOR4_X1 port map( A1 => n24973, A2 => n17484, A3 => n17471, A4 => 
                           n17472, ZN => n24974);
   U18302 : AND3_X1 port map( A1 => n24976, A2 => n24975, A3 => n24974, ZN => 
                           n24977);
   U18303 : OAI222_X1 port map( A1 => n19567, A2 => n22933, B1 => n24977, B2 =>
                           n22800, C1 => n19695, C2 => n22520, ZN => n24978);
   U18304 : AOI221_X1 port map( B1 => n22921, B2 => n22118, C1 => n22975, C2 =>
                           n21124, A => n24978, ZN => n24986);
   U18305 : OAI22_X1 port map( A1 => n19183, A2 => n22976, B1 => n19311, B2 => 
                           n22650, ZN => n24979);
   U18306 : OAI222_X1 port map( A1 => n18991, A2 => n22954, B1 => n19247, B2 =>
                           n22968, C1 => n19119, C2 => n22637, ZN => n24980);
   U18307 : AOI221_X1 port map( B1 => n22801, B2 => n22052, C1 => n22961, C2 =>
                           n21240, A => n24980, ZN => n24984);
   U18308 : OAI22_X1 port map( A1 => n23269, A2 => n24981, B1 => n18735, B2 => 
                           n22946, ZN => n24982);
   U18309 : AOI221_X1 port map( B1 => n23278, B2 => n20929, C1 => n22494, C2 =>
                           n21669, A => n24982, ZN => n24983);
   U18310 : NAND4_X1 port map( A1 => n24983, A2 => n24985, A3 => n24984, A4 => 
                           n24986, ZN => n3313);
   U18311 : NAND2_X1 port map( A1 => n17448, A2 => n17449, ZN => n24988);
   U18312 : AOI21_X1 port map( B1 => n17452, B2 => n17453, A => n23199, ZN => 
                           n24987);
   U18313 : AOI221_X1 port map( B1 => n23215, B2 => n21851, C1 => n23207, C2 =>
                           n24988, A => n24987, ZN => n24992);
   U18314 : AOI222_X1 port map( A1 => n23239, A2 => n21294, B1 => n23231, B2 =>
                           n20970, C1 => n23223, C2 => n20777, ZN => n24991);
   U18315 : OAI222_X1 port map( A1 => n20424, A2 => n23263, B1 => n20552, B2 =>
                           n23255, C1 => n20488, C2 => n23247, ZN => n24989);
   U18316 : NOR4_X1 port map( A1 => n24989, A2 => n17457, A3 => n17444, A4 => 
                           n17445, ZN => n24990);
   U18317 : AND3_X1 port map( A1 => n24992, A2 => n24991, A3 => n24990, ZN => 
                           n24993);
   U18318 : OAI222_X1 port map( A1 => n19528, A2 => n22937, B1 => n24993, B2 =>
                           n22798, C1 => n19656, C2 => n22518, ZN => n24994);
   U18319 : AOI221_X1 port map( B1 => n22921, B2 => n22119, C1 => n22970, C2 =>
                           n21101, A => n24994, ZN => n25002);
   U18320 : OAI22_X1 port map( A1 => n19144, A2 => n22980, B1 => n19272, B2 => 
                           n22640, ZN => n24995);
   U18321 : AOI221_X1 port map( B1 => n22920, B2 => n22076, C1 => n22803, C2 =>
                           n21155, A => n24995, ZN => n25001);
   U18322 : OAI222_X1 port map( A1 => n18952, A2 => n22954, B1 => n19208, B2 =>
                           n22964, C1 => n19080, C2 => n22635, ZN => n24996);
   U18323 : AOI221_X1 port map( B1 => n25391, B2 => n22165, C1 => n22962, C2 =>
                           n21217, A => n24996, ZN => n25000);
   U18324 : OAI22_X1 port map( A1 => n25394, A2 => n24997, B1 => n18696, B2 => 
                           n22946, ZN => n24998);
   U18325 : AOI221_X1 port map( B1 => n23278, B2 => n20906, C1 => n22494, C2 =>
                           n21646, A => n24998, ZN => n24999);
   U18326 : NAND4_X1 port map( A1 => n25000, A2 => n25001, A3 => n24999, A4 => 
                           n25002, ZN => n3314);
   U18327 : NAND2_X1 port map( A1 => n17421, A2 => n17422, ZN => n25004);
   U18328 : AOI21_X1 port map( B1 => n17425, B2 => n17426, A => n23199, ZN => 
                           n25003);
   U18329 : AOI221_X1 port map( B1 => n23215, B2 => n21903, C1 => n23207, C2 =>
                           n25004, A => n25003, ZN => n25008);
   U18330 : AOI222_X1 port map( A1 => n23239, A2 => n21346, B1 => n23231, B2 =>
                           n21022, C1 => n23223, C2 => n20829, ZN => n25007);
   U18331 : OAI222_X1 port map( A1 => n20464, A2 => n23263, B1 => n20592, B2 =>
                           n23255, C1 => n20528, C2 => n23247, ZN => n25005);
   U18332 : NOR4_X1 port map( A1 => n25005, A2 => n17430, A3 => n17417, A4 => 
                           n17418, ZN => n25006);
   U18333 : AND3_X1 port map( A1 => n25008, A2 => n25007, A3 => n25006, ZN => 
                           n25009);
   U18334 : OAI222_X1 port map( A1 => n19568, A2 => n22935, B1 => n25009, B2 =>
                           n22798, C1 => n19696, C2 => n22516, ZN => n25010);
   U18335 : OAI22_X1 port map( A1 => n19184, A2 => n22980, B1 => n19312, B2 => 
                           n22643, ZN => n25011);
   U18336 : AOI221_X1 port map( B1 => n22919, B2 => n22077, C1 => n22811, C2 =>
                           n21273, A => n25011, ZN => n25017);
   U18337 : OAI222_X1 port map( A1 => n18992, A2 => n22953, B1 => n19248, B2 =>
                           n22966, C1 => n19120, C2 => n22635, ZN => n25012);
   U18338 : AOI221_X1 port map( B1 => n25391, B2 => n22166, C1 => n22958, C2 =>
                           n21280, A => n25012, ZN => n25016);
   U18339 : OAI22_X1 port map( A1 => n23269, A2 => n25013, B1 => n18736, B2 => 
                           n22943, ZN => n25014);
   U18340 : AOI221_X1 port map( B1 => n23278, B2 => n20958, C1 => n22494, C2 =>
                           n21831, A => n25014, ZN => n25015);
   U18341 : NAND4_X1 port map( A1 => n25016, A2 => n25017, A3 => n25015, A4 => 
                           n25018, ZN => n3315);
   U18342 : NAND2_X1 port map( A1 => n17394, A2 => n17395, ZN => n25020);
   U18343 : AOI21_X1 port map( B1 => n17398, B2 => n17399, A => n23199, ZN => 
                           n25019);
   U18344 : AOI221_X1 port map( B1 => n23215, B2 => n21886, C1 => n23207, C2 =>
                           n25020, A => n25019, ZN => n25024);
   U18345 : AOI222_X1 port map( A1 => n23239, A2 => n21329, B1 => n23231, B2 =>
                           n21005, C1 => n23223, C2 => n20812, ZN => n25023);
   U18346 : OAI222_X1 port map( A1 => n20423, A2 => n23263, B1 => n20551, B2 =>
                           n23255, C1 => n20487, C2 => n23247, ZN => n25021);
   U18347 : NOR4_X1 port map( A1 => n25021, A2 => n17403, A3 => n17390, A4 => 
                           n17391, ZN => n25022);
   U18348 : AND3_X1 port map( A1 => n25024, A2 => n25023, A3 => n25022, ZN => 
                           n25025);
   U18349 : OAI222_X1 port map( A1 => n19527, A2 => n22935, B1 => n25025, B2 =>
                           n22799, C1 => n19655, C2 => n22521, ZN => n25026);
   U18350 : AOI221_X1 port map( B1 => n22923, B2 => n22120, C1 => n22975, C2 =>
                           n21135, A => n25026, ZN => n25034);
   U18351 : OAI22_X1 port map( A1 => n19143, A2 => n22976, B1 => n19271, B2 => 
                           n22632, ZN => n25027);
   U18352 : AOI221_X1 port map( B1 => n22914, B2 => n22078, C1 => n22807, C2 =>
                           n21169, A => n25027, ZN => n25033);
   U18353 : OAI222_X1 port map( A1 => n18951, A2 => n22954, B1 => n19207, B2 =>
                           n22964, C1 => n19079, C2 => n22636, ZN => n25028);
   U18354 : AOI221_X1 port map( B1 => n22801, B2 => n22053, C1 => n22962, C2 =>
                           n21253, A => n25028, ZN => n25032);
   U18355 : OAI22_X1 port map( A1 => n23269, A2 => n25029, B1 => n18695, B2 => 
                           n22944, ZN => n25030);
   U18356 : AOI221_X1 port map( B1 => n23278, B2 => n20941, C1 => n22494, C2 =>
                           n21681, A => n25030, ZN => n25031);
   U18357 : NAND4_X1 port map( A1 => n25031, A2 => n25033, A3 => n25032, A4 => 
                           n25034, ZN => n3316);
   U18358 : NAND2_X1 port map( A1 => n17367, A2 => n17368, ZN => n25036);
   U18359 : AOI21_X1 port map( B1 => n17371, B2 => n17372, A => n23199, ZN => 
                           n25035);
   U18360 : AOI221_X1 port map( B1 => n23215, B2 => n21852, C1 => n23207, C2 =>
                           n25036, A => n25035, ZN => n25040);
   U18361 : AOI222_X1 port map( A1 => n23239, A2 => n21295, B1 => n23231, B2 =>
                           n20971, C1 => n23223, C2 => n20778, ZN => n25039);
   U18362 : OAI222_X1 port map( A1 => n20465, A2 => n23263, B1 => n20593, B2 =>
                           n23255, C1 => n20529, C2 => n23247, ZN => n25037);
   U18363 : NOR4_X1 port map( A1 => n25037, A2 => n17376, A3 => n17363, A4 => 
                           n17364, ZN => n25038);
   U18364 : AND3_X1 port map( A1 => n25040, A2 => n25039, A3 => n25038, ZN => 
                           n25041);
   U18365 : OAI222_X1 port map( A1 => n19569, A2 => n22652, B1 => n25041, B2 =>
                           n22798, C1 => n19697, C2 => n22516, ZN => n25042);
   U18366 : AOI221_X1 port map( B1 => n22922, B2 => n22121, C1 => n22975, C2 =>
                           n21102, A => n25042, ZN => n25050);
   U18367 : OAI22_X1 port map( A1 => n19185, A2 => n22979, B1 => n19313, B2 => 
                           n22631, ZN => n25043);
   U18368 : AOI221_X1 port map( B1 => n22911, B2 => n22079, C1 => n22808, C2 =>
                           n21156, A => n25043, ZN => n25049);
   U18369 : OAI222_X1 port map( A1 => n18993, A2 => n22952, B1 => n19249, B2 =>
                           n22965, C1 => n19121, C2 => n22636, ZN => n25044);
   U18370 : AOI221_X1 port map( B1 => n25391, B2 => n22167, C1 => n22960, C2 =>
                           n21218, A => n25044, ZN => n25048);
   U18371 : OAI22_X1 port map( A1 => n23269, A2 => n25045, B1 => n18737, B2 => 
                           n22945, ZN => n25046);
   U18372 : AOI221_X1 port map( B1 => n23278, B2 => n20907, C1 => n22494, C2 =>
                           n21647, A => n25046, ZN => n25047);
   U18373 : NAND4_X1 port map( A1 => n25048, A2 => n25049, A3 => n25047, A4 => 
                           n25050, ZN => n3317);
   U18374 : NAND2_X1 port map( A1 => n17340, A2 => n17341, ZN => n25052);
   U18375 : AOI21_X1 port map( B1 => n17344, B2 => n17345, A => n23199, ZN => 
                           n25051);
   U18376 : AOI221_X1 port map( B1 => n23215, B2 => n21887, C1 => n23207, C2 =>
                           n25052, A => n25051, ZN => n25056);
   U18377 : AOI222_X1 port map( A1 => n23239, A2 => n21330, B1 => n23231, B2 =>
                           n21006, C1 => n23223, C2 => n20813, ZN => n25055);
   U18378 : OAI222_X1 port map( A1 => n20422, A2 => n23263, B1 => n20550, B2 =>
                           n23255, C1 => n20486, C2 => n23247, ZN => n25053);
   U18379 : NOR4_X1 port map( A1 => n25053, A2 => n17349, A3 => n17336, A4 => 
                           n17337, ZN => n25054);
   U18380 : AND3_X1 port map( A1 => n25056, A2 => n25055, A3 => n25054, ZN => 
                           n25057);
   U18381 : OAI222_X1 port map( A1 => n19526, A2 => n22933, B1 => n25057, B2 =>
                           n22799, C1 => n19654, C2 => n22519, ZN => n25058);
   U18382 : AOI221_X1 port map( B1 => n22523, B2 => n22122, C1 => n22975, C2 =>
                           n21136, A => n25058, ZN => n25066);
   U18383 : OAI22_X1 port map( A1 => n19142, A2 => n22978, B1 => n19270, B2 => 
                           n22630, ZN => n25059);
   U18384 : AOI221_X1 port map( B1 => n22920, B2 => n22080, C1 => n22807, C2 =>
                           n21170, A => n25059, ZN => n25065);
   U18385 : OAI222_X1 port map( A1 => n18950, A2 => n22953, B1 => n19206, B2 =>
                           n22966, C1 => n19078, C2 => n22636, ZN => n25060);
   U18386 : AOI221_X1 port map( B1 => n25391, B2 => n22168, C1 => n22961, C2 =>
                           n21254, A => n25060, ZN => n25064);
   U18387 : OAI22_X1 port map( A1 => n23269, A2 => n25061, B1 => n18694, B2 => 
                           n22946, ZN => n25062);
   U18388 : AOI221_X1 port map( B1 => n23278, B2 => n20942, C1 => n22494, C2 =>
                           n21682, A => n25062, ZN => n25063);
   U18389 : NAND4_X1 port map( A1 => n25064, A2 => n25065, A3 => n25063, A4 => 
                           n25066, ZN => n3318);
   U18390 : NAND2_X1 port map( A1 => n17313, A2 => n17314, ZN => n25068);
   U18391 : AOI21_X1 port map( B1 => n17317, B2 => n17318, A => n23199, ZN => 
                           n25067);
   U18392 : AOI221_X1 port map( B1 => n23215, B2 => n21853, C1 => n23207, C2 =>
                           n25068, A => n25067, ZN => n25072);
   U18393 : AOI222_X1 port map( A1 => n23239, A2 => n21296, B1 => n23231, B2 =>
                           n20972, C1 => n23223, C2 => n20779, ZN => n25071);
   U18394 : OAI222_X1 port map( A1 => n20466, A2 => n23263, B1 => n20594, B2 =>
                           n23255, C1 => n20530, C2 => n23247, ZN => n25069);
   U18395 : NOR4_X1 port map( A1 => n25069, A2 => n17322, A3 => n17309, A4 => 
                           n17310, ZN => n25070);
   U18396 : AND3_X1 port map( A1 => n25072, A2 => n25071, A3 => n25070, ZN => 
                           n25073);
   U18397 : OAI222_X1 port map( A1 => n19570, A2 => n22933, B1 => n25073, B2 =>
                           n22798, C1 => n19698, C2 => n22520, ZN => n25074);
   U18398 : AOI221_X1 port map( B1 => n22522, B2 => n22123, C1 => n22972, C2 =>
                           n21103, A => n25074, ZN => n25082);
   U18399 : OAI22_X1 port map( A1 => n19186, A2 => n22977, B1 => n19314, B2 => 
                           n22630, ZN => n25075);
   U18400 : AOI221_X1 port map( B1 => n22920, B2 => n22081, C1 => n22804, C2 =>
                           n21157, A => n25075, ZN => n25081);
   U18401 : OAI222_X1 port map( A1 => n18994, A2 => n22952, B1 => n19250, B2 =>
                           n22964, C1 => n19122, C2 => n22639, ZN => n25076);
   U18402 : AOI221_X1 port map( B1 => n25391, B2 => n22169, C1 => n22958, C2 =>
                           n21219, A => n25076, ZN => n25080);
   U18403 : OAI22_X1 port map( A1 => n23269, A2 => n25077, B1 => n18738, B2 => 
                           n22947, ZN => n25078);
   U18404 : AOI221_X1 port map( B1 => n23278, B2 => n20908, C1 => n22494, C2 =>
                           n21648, A => n25078, ZN => n25079);
   U18405 : NAND4_X1 port map( A1 => n25080, A2 => n25081, A3 => n25079, A4 => 
                           n25082, ZN => n3319);
   U18406 : NAND2_X1 port map( A1 => n17286, A2 => n17287, ZN => n25084);
   U18407 : AOI21_X1 port map( B1 => n17290, B2 => n17291, A => n23199, ZN => 
                           n25083);
   U18408 : AOI221_X1 port map( B1 => n23215, B2 => n21888, C1 => n23207, C2 =>
                           n25084, A => n25083, ZN => n25088);
   U18409 : AOI222_X1 port map( A1 => n23239, A2 => n21331, B1 => n23231, B2 =>
                           n21007, C1 => n23223, C2 => n20814, ZN => n25087);
   U18410 : OAI222_X1 port map( A1 => n20421, A2 => n23263, B1 => n20549, B2 =>
                           n23255, C1 => n20485, C2 => n23247, ZN => n25085);
   U18411 : NOR4_X1 port map( A1 => n25085, A2 => n17295, A3 => n17282, A4 => 
                           n17283, ZN => n25086);
   U18412 : AND3_X1 port map( A1 => n25088, A2 => n25087, A3 => n25086, ZN => 
                           n25089);
   U18413 : OAI222_X1 port map( A1 => n19525, A2 => n22934, B1 => n25089, B2 =>
                           n22799, C1 => n19653, C2 => n22516, ZN => n25090);
   U18414 : AOI221_X1 port map( B1 => n22923, B2 => n22124, C1 => n22970, C2 =>
                           n21137, A => n25090, ZN => n25098);
   U18415 : OAI22_X1 port map( A1 => n19141, A2 => n22979, B1 => n19269, B2 => 
                           n22648, ZN => n25091);
   U18416 : OAI222_X1 port map( A1 => n18949, A2 => n22951, B1 => n19205, B2 =>
                           n22964, C1 => n19077, C2 => n22637, ZN => n25092);
   U18417 : AOI221_X1 port map( B1 => n25391, B2 => n22170, C1 => n22962, C2 =>
                           n21255, A => n25092, ZN => n25096);
   U18418 : OAI22_X1 port map( A1 => n23269, A2 => n25093, B1 => n18693, B2 => 
                           n22944, ZN => n25094);
   U18419 : AOI221_X1 port map( B1 => n23278, B2 => n20943, C1 => n22494, C2 =>
                           n21683, A => n25094, ZN => n25095);
   U18420 : NAND4_X1 port map( A1 => n25096, A2 => n25097, A3 => n25095, A4 => 
                           n25098, ZN => n3320);
   U18421 : NAND2_X1 port map( A1 => n17259, A2 => n17260, ZN => n25100);
   U18422 : AOI21_X1 port map( B1 => n17263, B2 => n17264, A => n23199, ZN => 
                           n25099);
   U18423 : AOI221_X1 port map( B1 => n23215, B2 => n21889, C1 => n23207, C2 =>
                           n25100, A => n25099, ZN => n25104);
   U18424 : AOI222_X1 port map( A1 => n23239, A2 => n21332, B1 => n23231, B2 =>
                           n21008, C1 => n23223, C2 => n20815, ZN => n25103);
   U18425 : OAI222_X1 port map( A1 => n20467, A2 => n23263, B1 => n20595, B2 =>
                           n23255, C1 => n20531, C2 => n23247, ZN => n25101);
   U18426 : NOR4_X1 port map( A1 => n25101, A2 => n17268, A3 => n17255, A4 => 
                           n17256, ZN => n25102);
   U18427 : AND3_X1 port map( A1 => n25104, A2 => n25103, A3 => n25102, ZN => 
                           n25105);
   U18428 : OAI222_X1 port map( A1 => n19571, A2 => n22936, B1 => n25105, B2 =>
                           n22799, C1 => n19699, C2 => n22516, ZN => n25106);
   U18429 : AOI221_X1 port map( B1 => n22921, B2 => n22125, C1 => n22971, C2 =>
                           n21138, A => n25106, ZN => n25114);
   U18430 : OAI22_X1 port map( A1 => n19187, A2 => n22980, B1 => n19315, B2 => 
                           n22632, ZN => n25107);
   U18431 : AOI221_X1 port map( B1 => n22918, B2 => n22082, C1 => n22802, C2 =>
                           n21171, A => n25107, ZN => n25113);
   U18432 : OAI222_X1 port map( A1 => n18995, A2 => n22951, B1 => n19251, B2 =>
                           n22968, C1 => n19123, C2 => n22636, ZN => n25108);
   U18433 : AOI221_X1 port map( B1 => n25391, B2 => n22171, C1 => n22961, C2 =>
                           n21256, A => n25108, ZN => n25112);
   U18434 : OAI22_X1 port map( A1 => n23269, A2 => n25109, B1 => n18739, B2 => 
                           n22945, ZN => n25110);
   U18435 : AOI221_X1 port map( B1 => n23278, B2 => n20944, C1 => n22494, C2 =>
                           n21684, A => n25110, ZN => n25111);
   U18436 : NAND4_X1 port map( A1 => n25112, A2 => n25113, A3 => n25111, A4 => 
                           n25114, ZN => n3321);
   U18437 : NAND2_X1 port map( A1 => n17232, A2 => n17233, ZN => n25116);
   U18438 : AOI21_X1 port map( B1 => n17236, B2 => n17237, A => n23199, ZN => 
                           n25115);
   U18439 : AOI221_X1 port map( B1 => n23215, B2 => n21854, C1 => n23207, C2 =>
                           n25116, A => n25115, ZN => n25120);
   U18440 : AOI222_X1 port map( A1 => n23239, A2 => n21297, B1 => n23231, B2 =>
                           n20973, C1 => n23223, C2 => n20780, ZN => n25119);
   U18441 : OAI222_X1 port map( A1 => n20420, A2 => n23263, B1 => n20548, B2 =>
                           n23255, C1 => n20484, C2 => n23247, ZN => n25117);
   U18442 : NOR4_X1 port map( A1 => n25117, A2 => n17241, A3 => n17228, A4 => 
                           n17229, ZN => n25118);
   U18443 : AND3_X1 port map( A1 => n25120, A2 => n25119, A3 => n25118, ZN => 
                           n25121);
   U18444 : OAI222_X1 port map( A1 => n19524, A2 => n22652, B1 => n25121, B2 =>
                           n22798, C1 => n19652, C2 => n22519, ZN => n25122);
   U18445 : AOI221_X1 port map( B1 => n22922, B2 => n22126, C1 => n22972, C2 =>
                           n21104, A => n25122, ZN => n25130);
   U18446 : OAI22_X1 port map( A1 => n19140, A2 => n22976, B1 => n19268, B2 => 
                           n22633, ZN => n25123);
   U18447 : OAI222_X1 port map( A1 => n18948, A2 => n22952, B1 => n19204, B2 =>
                           n22964, C1 => n19076, C2 => n22636, ZN => n25124);
   U18448 : AOI221_X1 port map( B1 => n25391, B2 => n22172, C1 => n22962, C2 =>
                           n21220, A => n25124, ZN => n25128);
   U18449 : OAI22_X1 port map( A1 => n23269, A2 => n25125, B1 => n18692, B2 => 
                           n22943, ZN => n25126);
   U18450 : AOI221_X1 port map( B1 => n23278, B2 => n20909, C1 => n22494, C2 =>
                           n21649, A => n25126, ZN => n25127);
   U18451 : NAND4_X1 port map( A1 => n25128, A2 => n25129, A3 => n25127, A4 => 
                           n25130, ZN => n3322);
   U18452 : NAND2_X1 port map( A1 => n17205, A2 => n17206, ZN => n25132);
   U18453 : AOI21_X1 port map( B1 => n17209, B2 => n17210, A => n23200, ZN => 
                           n25131);
   U18454 : AOI221_X1 port map( B1 => n23216, B2 => n21890, C1 => n23208, C2 =>
                           n25132, A => n25131, ZN => n25136);
   U18455 : AOI222_X1 port map( A1 => n23240, A2 => n21333, B1 => n23232, B2 =>
                           n21009, C1 => n23224, C2 => n20816, ZN => n25135);
   U18456 : OAI222_X1 port map( A1 => n20468, A2 => n23264, B1 => n20596, B2 =>
                           n23256, C1 => n20532, C2 => n23248, ZN => n25133);
   U18457 : NOR4_X1 port map( A1 => n25133, A2 => n17214, A3 => n17201, A4 => 
                           n17202, ZN => n25134);
   U18458 : AND3_X1 port map( A1 => n25136, A2 => n25135, A3 => n25134, ZN => 
                           n25137);
   U18459 : OAI222_X1 port map( A1 => n19572, A2 => n22933, B1 => n25137, B2 =>
                           n22799, C1 => n19700, C2 => n22516, ZN => n25138);
   U18460 : AOI221_X1 port map( B1 => n22523, B2 => n22127, C1 => n22973, C2 =>
                           n21139, A => n25138, ZN => n25146);
   U18461 : OAI22_X1 port map( A1 => n19188, A2 => n22980, B1 => n19316, B2 => 
                           n22629, ZN => n25139);
   U18462 : AOI221_X1 port map( B1 => n22918, B2 => n22083, C1 => n22811, C2 =>
                           n21172, A => n25139, ZN => n25145);
   U18463 : OAI222_X1 port map( A1 => n18996, A2 => n22951, B1 => n19252, B2 =>
                           n22965, C1 => n19124, C2 => n22637, ZN => n25140);
   U18464 : AOI221_X1 port map( B1 => n22801, B2 => n22054, C1 => n22957, C2 =>
                           n21257, A => n25140, ZN => n25144);
   U18465 : OAI22_X1 port map( A1 => n23269, A2 => n25141, B1 => n18740, B2 => 
                           n22944, ZN => n25142);
   U18466 : AOI221_X1 port map( B1 => n23279, B2 => n20945, C1 => n22494, C2 =>
                           n21685, A => n25142, ZN => n25143);
   U18467 : NAND4_X1 port map( A1 => n25143, A2 => n25145, A3 => n25144, A4 => 
                           n25146, ZN => n3323);
   U18468 : NAND2_X1 port map( A1 => n17178, A2 => n17179, ZN => n25148);
   U18469 : AOI21_X1 port map( B1 => n17182, B2 => n17183, A => n23200, ZN => 
                           n25147);
   U18470 : AOI221_X1 port map( B1 => n23216, B2 => n21875, C1 => n23208, C2 =>
                           n25148, A => n25147, ZN => n25152);
   U18471 : AOI222_X1 port map( A1 => n23240, A2 => n21318, B1 => n23232, B2 =>
                           n20994, C1 => n23224, C2 => n20801, ZN => n25151);
   U18472 : OAI222_X1 port map( A1 => n20419, A2 => n23264, B1 => n20547, B2 =>
                           n23256, C1 => n20483, C2 => n23248, ZN => n25149);
   U18473 : NOR4_X1 port map( A1 => n25149, A2 => n17187, A3 => n17174, A4 => 
                           n17175, ZN => n25150);
   U18474 : AND3_X1 port map( A1 => n25152, A2 => n25151, A3 => n25150, ZN => 
                           n25153);
   U18475 : OAI222_X1 port map( A1 => n19523, A2 => n22935, B1 => n25153, B2 =>
                           n22800, C1 => n19651, C2 => n22517, ZN => n25154);
   U18476 : AOI221_X1 port map( B1 => n22522, B2 => n22128, C1 => n22974, C2 =>
                           n21125, A => n25154, ZN => n25162);
   U18477 : OAI22_X1 port map( A1 => n19139, A2 => n22979, B1 => n19267, B2 => 
                           n22648, ZN => n25155);
   U18478 : OAI222_X1 port map( A1 => n18947, A2 => n22954, B1 => n19203, B2 =>
                           n22965, C1 => n19075, C2 => n22638, ZN => n25156);
   U18479 : AOI221_X1 port map( B1 => n25391, B2 => n22173, C1 => n22957, C2 =>
                           n21241, A => n25156, ZN => n25160);
   U18480 : OAI22_X1 port map( A1 => n23269, A2 => n25157, B1 => n18691, B2 => 
                           n22945, ZN => n25158);
   U18481 : AOI221_X1 port map( B1 => n23279, B2 => n20930, C1 => n22494, C2 =>
                           n21670, A => n25158, ZN => n25159);
   U18482 : NAND4_X1 port map( A1 => n25160, A2 => n25161, A3 => n25159, A4 => 
                           n25162, ZN => n3324);
   U18483 : NAND2_X1 port map( A1 => n17151, A2 => n17152, ZN => n25164);
   U18484 : AOI21_X1 port map( B1 => n17155, B2 => n17156, A => n23200, ZN => 
                           n25163);
   U18485 : AOI221_X1 port map( B1 => n23216, B2 => n21855, C1 => n23208, C2 =>
                           n25164, A => n25163, ZN => n25168);
   U18486 : AOI222_X1 port map( A1 => n23240, A2 => n21298, B1 => n23232, B2 =>
                           n20974, C1 => n23224, C2 => n20781, ZN => n25167);
   U18487 : OAI222_X1 port map( A1 => n20469, A2 => n23264, B1 => n20597, B2 =>
                           n23256, C1 => n20533, C2 => n23248, ZN => n25165);
   U18488 : NOR4_X1 port map( A1 => n25165, A2 => n17160, A3 => n17147, A4 => 
                           n17148, ZN => n25166);
   U18489 : AND3_X1 port map( A1 => n25168, A2 => n25167, A3 => n25166, ZN => 
                           n25169);
   U18490 : OAI222_X1 port map( A1 => n19573, A2 => n22936, B1 => n25169, B2 =>
                           n22798, C1 => n19701, C2 => n22521, ZN => n25170);
   U18491 : AOI221_X1 port map( B1 => n22522, B2 => n22129, C1 => n22975, C2 =>
                           n21105, A => n25170, ZN => n25178);
   U18492 : OAI22_X1 port map( A1 => n19189, A2 => n22978, B1 => n19317, B2 => 
                           n22650, ZN => n25171);
   U18493 : OAI222_X1 port map( A1 => n18997, A2 => n22954, B1 => n19253, B2 =>
                           n22967, C1 => n19125, C2 => n22635, ZN => n25172);
   U18494 : AOI221_X1 port map( B1 => n25391, B2 => n22174, C1 => n22958, C2 =>
                           n21221, A => n25172, ZN => n25176);
   U18495 : OAI22_X1 port map( A1 => n23269, A2 => n25173, B1 => n18741, B2 => 
                           n22945, ZN => n25174);
   U18496 : AOI221_X1 port map( B1 => n23279, B2 => n20910, C1 => n22494, C2 =>
                           n21650, A => n25174, ZN => n25175);
   U18497 : NAND4_X1 port map( A1 => n25176, A2 => n25177, A3 => n25175, A4 => 
                           n25178, ZN => n3325);
   U18498 : NAND2_X1 port map( A1 => n17124, A2 => n17125, ZN => n25180);
   U18499 : AOI21_X1 port map( B1 => n17128, B2 => n17129, A => n23200, ZN => 
                           n25179);
   U18500 : AOI221_X1 port map( B1 => n23216, B2 => n21891, C1 => n23208, C2 =>
                           n25180, A => n25179, ZN => n25184);
   U18501 : AOI222_X1 port map( A1 => n23240, A2 => n21334, B1 => n23232, B2 =>
                           n21010, C1 => n23224, C2 => n20817, ZN => n25183);
   U18502 : OAI222_X1 port map( A1 => n20418, A2 => n23264, B1 => n20546, B2 =>
                           n23256, C1 => n20482, C2 => n23248, ZN => n25181);
   U18503 : NOR4_X1 port map( A1 => n25181, A2 => n17133, A3 => n17120, A4 => 
                           n17121, ZN => n25182);
   U18504 : AND3_X1 port map( A1 => n25184, A2 => n25183, A3 => n25182, ZN => 
                           n25185);
   U18505 : OAI222_X1 port map( A1 => n19522, A2 => n22935, B1 => n25185, B2 =>
                           n22799, C1 => n19650, C2 => n22518, ZN => n25186);
   U18506 : AOI221_X1 port map( B1 => n22921, B2 => n22130, C1 => n22975, C2 =>
                           n21140, A => n25186, ZN => n25194);
   U18507 : OAI22_X1 port map( A1 => n19138, A2 => n22979, B1 => n19266, B2 => 
                           n22644, ZN => n25187);
   U18508 : OAI222_X1 port map( A1 => n18946, A2 => n22953, B1 => n19202, B2 =>
                           n22966, C1 => n19074, C2 => n22639, ZN => n25188);
   U18509 : AOI221_X1 port map( B1 => n25391, B2 => n22175, C1 => n22959, C2 =>
                           n21258, A => n25188, ZN => n25192);
   U18510 : OAI22_X1 port map( A1 => n23269, A2 => n25189, B1 => n18690, B2 => 
                           n22946, ZN => n25190);
   U18511 : AOI221_X1 port map( B1 => n23279, B2 => n20946, C1 => n22494, C2 =>
                           n21686, A => n25190, ZN => n25191);
   U18512 : NAND4_X1 port map( A1 => n25192, A2 => n25193, A3 => n25191, A4 => 
                           n25194, ZN => n3326);
   U18513 : NAND2_X1 port map( A1 => n17097, A2 => n17098, ZN => n25196);
   U18514 : AOI21_X1 port map( B1 => n17101, B2 => n17102, A => n23200, ZN => 
                           n25195);
   U18515 : AOI221_X1 port map( B1 => n23216, B2 => n21892, C1 => n23208, C2 =>
                           n25196, A => n25195, ZN => n25200);
   U18516 : AOI222_X1 port map( A1 => n23240, A2 => n21335, B1 => n23232, B2 =>
                           n21011, C1 => n23224, C2 => n20818, ZN => n25199);
   U18517 : OAI222_X1 port map( A1 => n20470, A2 => n23264, B1 => n20598, B2 =>
                           n23256, C1 => n20534, C2 => n23248, ZN => n25197);
   U18518 : NOR4_X1 port map( A1 => n25197, A2 => n17106, A3 => n17093, A4 => 
                           n17094, ZN => n25198);
   U18519 : AND3_X1 port map( A1 => n25200, A2 => n25199, A3 => n25198, ZN => 
                           n25201);
   U18520 : OAI222_X1 port map( A1 => n19574, A2 => n22936, B1 => n25201, B2 =>
                           n22799, C1 => n19702, C2 => n22517, ZN => n25202);
   U18521 : AOI221_X1 port map( B1 => n22921, B2 => n22131, C1 => n22975, C2 =>
                           n21141, A => n25202, ZN => n25210);
   U18522 : OAI22_X1 port map( A1 => n19190, A2 => n22978, B1 => n19318, B2 => 
                           n22641, ZN => n25203);
   U18523 : OAI222_X1 port map( A1 => n18998, A2 => n22952, B1 => n19254, B2 =>
                           n22965, C1 => n19126, C2 => n22638, ZN => n25204);
   U18524 : AOI221_X1 port map( B1 => n25391, B2 => n22176, C1 => n22960, C2 =>
                           n21259, A => n25204, ZN => n25208);
   U18525 : OAI22_X1 port map( A1 => n25394, A2 => n25205, B1 => n18742, B2 => 
                           n22947, ZN => n25206);
   U18526 : AOI221_X1 port map( B1 => n23279, B2 => n20947, C1 => n22494, C2 =>
                           n21687, A => n25206, ZN => n25207);
   U18527 : NAND4_X1 port map( A1 => n25208, A2 => n25209, A3 => n25207, A4 => 
                           n25210, ZN => n3327);
   U18528 : NAND2_X1 port map( A1 => n17070, A2 => n17071, ZN => n25212);
   U18529 : AOI21_X1 port map( B1 => n17074, B2 => n17075, A => n23200, ZN => 
                           n25211);
   U18530 : AOI221_X1 port map( B1 => n23216, B2 => n21856, C1 => n23208, C2 =>
                           n25212, A => n25211, ZN => n25216);
   U18531 : AOI222_X1 port map( A1 => n23240, A2 => n21299, B1 => n23232, B2 =>
                           n20975, C1 => n23224, C2 => n20782, ZN => n25215);
   U18532 : OAI222_X1 port map( A1 => n20417, A2 => n23264, B1 => n20545, B2 =>
                           n23256, C1 => n20481, C2 => n23248, ZN => n25213);
   U18533 : NOR4_X1 port map( A1 => n25213, A2 => n17079, A3 => n17066, A4 => 
                           n17067, ZN => n25214);
   U18534 : AND3_X1 port map( A1 => n25216, A2 => n25215, A3 => n25214, ZN => 
                           n25217);
   U18535 : OAI222_X1 port map( A1 => n19521, A2 => n22934, B1 => n25217, B2 =>
                           n22798, C1 => n19649, C2 => n22518, ZN => n25218);
   U18536 : AOI221_X1 port map( B1 => n22523, B2 => n22132, C1 => n22970, C2 =>
                           n21106, A => n25218, ZN => n25226);
   U18537 : OAI22_X1 port map( A1 => n19137, A2 => n22977, B1 => n19265, B2 => 
                           n22645, ZN => n25219);
   U18538 : OAI222_X1 port map( A1 => n18945, A2 => n22955, B1 => n19201, B2 =>
                           n22966, C1 => n19073, C2 => n22636, ZN => n25220);
   U18539 : AOI221_X1 port map( B1 => n22801, B2 => n22055, C1 => n22961, C2 =>
                           n21222, A => n25220, ZN => n25224);
   U18540 : OAI22_X1 port map( A1 => n23270, A2 => n25221, B1 => n18689, B2 => 
                           n22943, ZN => n25222);
   U18541 : AOI221_X1 port map( B1 => n23279, B2 => n20911, C1 => n22494, C2 =>
                           n21651, A => n25222, ZN => n25223);
   U18542 : NAND4_X1 port map( A1 => n25223, A2 => n25225, A3 => n25224, A4 => 
                           n25226, ZN => n3328);
   U18543 : NAND2_X1 port map( A1 => n17043, A2 => n17044, ZN => n25228);
   U18544 : AOI21_X1 port map( B1 => n17047, B2 => n17048, A => n23200, ZN => 
                           n25227);
   U18545 : AOI221_X1 port map( B1 => n23216, B2 => n21893, C1 => n23208, C2 =>
                           n25228, A => n25227, ZN => n25232);
   U18546 : AOI222_X1 port map( A1 => n23240, A2 => n21336, B1 => n23232, B2 =>
                           n21012, C1 => n23224, C2 => n20819, ZN => n25231);
   U18547 : OAI222_X1 port map( A1 => n20471, A2 => n23264, B1 => n20599, B2 =>
                           n23256, C1 => n20535, C2 => n23248, ZN => n25229);
   U18548 : NOR4_X1 port map( A1 => n25229, A2 => n17052, A3 => n17039, A4 => 
                           n17040, ZN => n25230);
   U18549 : AND3_X1 port map( A1 => n25232, A2 => n25231, A3 => n25230, ZN => 
                           n25233);
   U18550 : OAI222_X1 port map( A1 => n19575, A2 => n22937, B1 => n25233, B2 =>
                           n22799, C1 => n19703, C2 => n22516, ZN => n25234);
   U18551 : AOI221_X1 port map( B1 => n22923, B2 => n22133, C1 => n22973, C2 =>
                           n21142, A => n25234, ZN => n25242);
   U18552 : OAI22_X1 port map( A1 => n19191, A2 => n22976, B1 => n19319, B2 => 
                           n22651, ZN => n25235);
   U18553 : OAI222_X1 port map( A1 => n18999, A2 => n22953, B1 => n19255, B2 =>
                           n22966, C1 => n19127, C2 => n22638, ZN => n25236);
   U18554 : AOI221_X1 port map( B1 => n25391, B2 => n22177, C1 => n22961, C2 =>
                           n21260, A => n25236, ZN => n25240);
   U18555 : OAI22_X1 port map( A1 => n25394, A2 => n25237, B1 => n18743, B2 => 
                           n22946, ZN => n25238);
   U18556 : AOI221_X1 port map( B1 => n23279, B2 => n20948, C1 => n22494, C2 =>
                           n21688, A => n25238, ZN => n25239);
   U18557 : NAND4_X1 port map( A1 => n25240, A2 => n25241, A3 => n25239, A4 => 
                           n25242, ZN => n3329);
   U18558 : NAND2_X1 port map( A1 => n17016, A2 => n17017, ZN => n25244);
   U18559 : AOI21_X1 port map( B1 => n17020, B2 => n17021, A => n23200, ZN => 
                           n25243);
   U18560 : AOI221_X1 port map( B1 => n23216, B2 => n21894, C1 => n23208, C2 =>
                           n25244, A => n25243, ZN => n25248);
   U18561 : AOI222_X1 port map( A1 => n23240, A2 => n21337, B1 => n23232, B2 =>
                           n21013, C1 => n23224, C2 => n20820, ZN => n25247);
   U18562 : OAI222_X1 port map( A1 => n20416, A2 => n23264, B1 => n20544, B2 =>
                           n23256, C1 => n20480, C2 => n23248, ZN => n25245);
   U18563 : NOR4_X1 port map( A1 => n25245, A2 => n17025, A3 => n17012, A4 => 
                           n17013, ZN => n25246);
   U18564 : AND3_X1 port map( A1 => n25248, A2 => n25247, A3 => n25246, ZN => 
                           n25249);
   U18565 : OAI222_X1 port map( A1 => n19520, A2 => n22935, B1 => n25249, B2 =>
                           n22799, C1 => n19648, C2 => n22520, ZN => n25250);
   U18566 : AOI221_X1 port map( B1 => n22923, B2 => n22134, C1 => n22972, C2 =>
                           n21143, A => n25250, ZN => n25258);
   U18567 : OAI22_X1 port map( A1 => n19136, A2 => n22977, B1 => n19264, B2 => 
                           n22645, ZN => n25251);
   U18568 : OAI222_X1 port map( A1 => n18944, A2 => n22953, B1 => n19200, B2 =>
                           n22966, C1 => n19072, C2 => n22638, ZN => n25252);
   U18569 : OAI22_X1 port map( A1 => n23270, A2 => n25253, B1 => n18688, B2 => 
                           n22947, ZN => n25254);
   U18570 : AOI221_X1 port map( B1 => n23279, B2 => n20949, C1 => n22494, C2 =>
                           n21689, A => n25254, ZN => n25255);
   U18571 : NAND4_X1 port map( A1 => n25255, A2 => n25257, A3 => n25256, A4 => 
                           n25258, ZN => n3330);
   U18572 : NAND2_X1 port map( A1 => n16989, A2 => n16990, ZN => n25260);
   U18573 : AOI21_X1 port map( B1 => n16993, B2 => n16994, A => n23200, ZN => 
                           n25259);
   U18574 : AOI221_X1 port map( B1 => n23216, B2 => n21857, C1 => n23208, C2 =>
                           n25260, A => n25259, ZN => n25264);
   U18575 : AOI222_X1 port map( A1 => n23240, A2 => n21300, B1 => n23232, B2 =>
                           n20976, C1 => n23224, C2 => n20783, ZN => n25263);
   U18576 : OAI222_X1 port map( A1 => n20472, A2 => n23264, B1 => n20600, B2 =>
                           n23256, C1 => n20536, C2 => n23248, ZN => n25261);
   U18577 : NOR4_X1 port map( A1 => n25261, A2 => n16998, A3 => n16985, A4 => 
                           n16986, ZN => n25262);
   U18578 : AND3_X1 port map( A1 => n25264, A2 => n25263, A3 => n25262, ZN => 
                           n25265);
   U18579 : OAI222_X1 port map( A1 => n19576, A2 => n22933, B1 => n25265, B2 =>
                           n22798, C1 => n19704, C2 => n22517, ZN => n25266);
   U18580 : AOI221_X1 port map( B1 => n22922, B2 => n22135, C1 => n22975, C2 =>
                           n21107, A => n25266, ZN => n25274);
   U18581 : OAI22_X1 port map( A1 => n19192, A2 => n22978, B1 => n19320, B2 => 
                           n22645, ZN => n25267);
   U18582 : OAI222_X1 port map( A1 => n19000, A2 => n22951, B1 => n19256, B2 =>
                           n22965, C1 => n19128, C2 => n22638, ZN => n25268);
   U18583 : AOI221_X1 port map( B1 => n25391, B2 => n22178, C1 => n22960, C2 =>
                           n21223, A => n25268, ZN => n25272);
   U18584 : OAI22_X1 port map( A1 => n25394, A2 => n25269, B1 => n18744, B2 => 
                           n22944, ZN => n25270);
   U18585 : AOI221_X1 port map( B1 => n23279, B2 => n20912, C1 => n22494, C2 =>
                           n21652, A => n25270, ZN => n25271);
   U18586 : NAND4_X1 port map( A1 => n25272, A2 => n25273, A3 => n25271, A4 => 
                           n25274, ZN => n3331);
   U18587 : NAND2_X1 port map( A1 => n16962, A2 => n16963, ZN => n25276);
   U18588 : AOI21_X1 port map( B1 => n16966, B2 => n16967, A => n23200, ZN => 
                           n25275);
   U18589 : AOI221_X1 port map( B1 => n23216, B2 => n21895, C1 => n23208, C2 =>
                           n25276, A => n25275, ZN => n25280);
   U18590 : AOI222_X1 port map( A1 => n23240, A2 => n21338, B1 => n23232, B2 =>
                           n21014, C1 => n23224, C2 => n20821, ZN => n25279);
   U18591 : OAI222_X1 port map( A1 => n20415, A2 => n23264, B1 => n20543, B2 =>
                           n23256, C1 => n20479, C2 => n23248, ZN => n25277);
   U18592 : NOR4_X1 port map( A1 => n25277, A2 => n16971, A3 => n16958, A4 => 
                           n16959, ZN => n25278);
   U18593 : AND3_X1 port map( A1 => n25280, A2 => n25279, A3 => n25278, ZN => 
                           n25281);
   U18594 : OAI222_X1 port map( A1 => n19519, A2 => n22652, B1 => n25281, B2 =>
                           n22799, C1 => n19647, C2 => n22521, ZN => n25282);
   U18595 : AOI221_X1 port map( B1 => n22922, B2 => n22136, C1 => n22975, C2 =>
                           n21144, A => n25282, ZN => n25290);
   U18596 : OAI22_X1 port map( A1 => n19135, A2 => n22980, B1 => n19263, B2 => 
                           n22649, ZN => n25283);
   U18597 : AOI221_X1 port map( B1 => n22917, B2 => n22084, C1 => n22810, C2 =>
                           n21173, A => n25283, ZN => n25289);
   U18598 : OAI222_X1 port map( A1 => n18943, A2 => n22951, B1 => n19199, B2 =>
                           n22968, C1 => n19071, C2 => n22635, ZN => n25284);
   U18599 : AOI221_X1 port map( B1 => n25391, B2 => n22179, C1 => n22961, C2 =>
                           n21261, A => n25284, ZN => n25288);
   U18600 : OAI22_X1 port map( A1 => n25394, A2 => n25285, B1 => n18687, B2 => 
                           n22945, ZN => n25286);
   U18601 : AOI221_X1 port map( B1 => n23279, B2 => n20950, C1 => n22494, C2 =>
                           n21690, A => n25286, ZN => n25287);
   U18602 : NAND4_X1 port map( A1 => n25288, A2 => n25289, A3 => n25287, A4 => 
                           n25290, ZN => n3332);
   U18603 : NAND2_X1 port map( A1 => n16935, A2 => n16936, ZN => n25292);
   U18604 : AOI21_X1 port map( B1 => n16939, B2 => n16940, A => n23200, ZN => 
                           n25291);
   U18605 : AOI221_X1 port map( B1 => n23216, B2 => n21896, C1 => n23208, C2 =>
                           n25292, A => n25291, ZN => n25296);
   U18606 : AOI222_X1 port map( A1 => n23240, A2 => n21339, B1 => n23232, B2 =>
                           n21015, C1 => n23224, C2 => n20822, ZN => n25295);
   U18607 : OAI222_X1 port map( A1 => n20473, A2 => n23264, B1 => n20601, B2 =>
                           n23256, C1 => n20537, C2 => n23248, ZN => n25293);
   U18608 : NOR4_X1 port map( A1 => n25293, A2 => n16944, A3 => n16931, A4 => 
                           n16932, ZN => n25294);
   U18609 : AND3_X1 port map( A1 => n25296, A2 => n25295, A3 => n25294, ZN => 
                           n25297);
   U18610 : OAI222_X1 port map( A1 => n19577, A2 => n22936, B1 => n25297, B2 =>
                           n22799, C1 => n19705, C2 => n22521, ZN => n25298);
   U18611 : AOI221_X1 port map( B1 => n22921, B2 => n22137, C1 => n22974, C2 =>
                           n21145, A => n25298, ZN => n25306);
   U18612 : OAI22_X1 port map( A1 => n19193, A2 => n22979, B1 => n19321, B2 => 
                           n22642, ZN => n25299);
   U18613 : OAI222_X1 port map( A1 => n19001, A2 => n22955, B1 => n19257, B2 =>
                           n22966, C1 => n19129, C2 => n22639, ZN => n25300);
   U18614 : AOI221_X1 port map( B1 => n25391, B2 => n22180, C1 => n22958, C2 =>
                           n21262, A => n25300, ZN => n25304);
   U18615 : OAI22_X1 port map( A1 => n25394, A2 => n25301, B1 => n18745, B2 => 
                           n22946, ZN => n25302);
   U18616 : AOI221_X1 port map( B1 => n23279, B2 => n20951, C1 => n22494, C2 =>
                           n21691, A => n25302, ZN => n25303);
   U18617 : NAND4_X1 port map( A1 => n25304, A2 => n25305, A3 => n25303, A4 => 
                           n25306, ZN => n3333);
   U18618 : NAND2_X1 port map( A1 => n16908, A2 => n16909, ZN => n25308);
   U18619 : AOI21_X1 port map( B1 => n16912, B2 => n16913, A => n23200, ZN => 
                           n25307);
   U18620 : AOI221_X1 port map( B1 => n23216, B2 => n21858, C1 => n23208, C2 =>
                           n25308, A => n25307, ZN => n25312);
   U18621 : AOI222_X1 port map( A1 => n23240, A2 => n21301, B1 => n23232, B2 =>
                           n20977, C1 => n23224, C2 => n20784, ZN => n25311);
   U18622 : OAI222_X1 port map( A1 => n20414, A2 => n23264, B1 => n20542, B2 =>
                           n23256, C1 => n20478, C2 => n23248, ZN => n25309);
   U18623 : NOR4_X1 port map( A1 => n25309, A2 => n16917, A3 => n16904, A4 => 
                           n16905, ZN => n25310);
   U18624 : AND3_X1 port map( A1 => n25312, A2 => n25311, A3 => n25310, ZN => 
                           n25313);
   U18625 : OAI222_X1 port map( A1 => n19518, A2 => n22934, B1 => n25313, B2 =>
                           n22798, C1 => n19646, C2 => n22520, ZN => n25314);
   U18626 : AOI221_X1 port map( B1 => n22923, B2 => n22138, C1 => n22975, C2 =>
                           n21108, A => n25314, ZN => n25322);
   U18627 : OAI22_X1 port map( A1 => n19134, A2 => n22978, B1 => n19262, B2 => 
                           n22651, ZN => n25315);
   U18628 : OAI222_X1 port map( A1 => n18942, A2 => n22954, B1 => n19198, B2 =>
                           n22965, C1 => n19070, C2 => n22635, ZN => n25316);
   U18629 : AOI221_X1 port map( B1 => n22801, B2 => n22056, C1 => n22962, C2 =>
                           n21224, A => n25316, ZN => n25320);
   U18630 : OAI22_X1 port map( A1 => n23270, A2 => n25317, B1 => n18686, B2 => 
                           n22947, ZN => n25318);
   U18631 : AOI221_X1 port map( B1 => n23279, B2 => n20913, C1 => n22494, C2 =>
                           n21653, A => n25318, ZN => n25319);
   U18632 : NAND4_X1 port map( A1 => n25319, A2 => n25321, A3 => n25320, A4 => 
                           n25322, ZN => n3334);
   U18633 : NAND2_X1 port map( A1 => n16881, A2 => n16882, ZN => n25324);
   U18634 : AOI21_X1 port map( B1 => n16885, B2 => n16886, A => n23201, ZN => 
                           n25323);
   U18635 : AOI221_X1 port map( B1 => n23217, B2 => n21897, C1 => n23209, C2 =>
                           n25324, A => n25323, ZN => n25328);
   U18636 : AOI222_X1 port map( A1 => n23241, A2 => n21340, B1 => n23233, B2 =>
                           n21016, C1 => n23225, C2 => n20823, ZN => n25327);
   U18637 : OAI222_X1 port map( A1 => n20474, A2 => n23265, B1 => n20602, B2 =>
                           n23257, C1 => n20538, C2 => n23249, ZN => n25325);
   U18638 : NOR4_X1 port map( A1 => n25325, A2 => n16890, A3 => n16877, A4 => 
                           n16878, ZN => n25326);
   U18639 : AND3_X1 port map( A1 => n25328, A2 => n25327, A3 => n25326, ZN => 
                           n25329);
   U18640 : OAI222_X1 port map( A1 => n19578, A2 => n22933, B1 => n25329, B2 =>
                           n22799, C1 => n19706, C2 => n22521, ZN => n25330);
   U18641 : AOI221_X1 port map( B1 => n22523, B2 => n22139, C1 => n22973, C2 =>
                           n21147, A => n25330, ZN => n25338);
   U18642 : OAI22_X1 port map( A1 => n19194, A2 => n22977, B1 => n19322, B2 => 
                           n22642, ZN => n25331);
   U18643 : OAI222_X1 port map( A1 => n19002, A2 => n22952, B1 => n19258, B2 =>
                           n22967, C1 => n19130, C2 => n22639, ZN => n25332);
   U18644 : AOI221_X1 port map( B1 => n25391, B2 => n22181, C1 => n22962, C2 =>
                           n21263, A => n25332, ZN => n25336);
   U18645 : OAI22_X1 port map( A1 => n25394, A2 => n25333, B1 => n18746, B2 => 
                           n22943, ZN => n25334);
   U18646 : AOI221_X1 port map( B1 => n23280, B2 => n20952, C1 => n22494, C2 =>
                           n21692, A => n25334, ZN => n25335);
   U18647 : NAND4_X1 port map( A1 => n25336, A2 => n25337, A3 => n25335, A4 => 
                           n25338, ZN => n3335);
   U18648 : NAND2_X1 port map( A1 => n16854, A2 => n16855, ZN => n25340);
   U18649 : AOI21_X1 port map( B1 => n16858, B2 => n16859, A => n23201, ZN => 
                           n25339);
   U18650 : AOI221_X1 port map( B1 => n23217, B2 => n21898, C1 => n23209, C2 =>
                           n25340, A => n25339, ZN => n25344);
   U18651 : AOI222_X1 port map( A1 => n23241, A2 => n21341, B1 => n23233, B2 =>
                           n21017, C1 => n23225, C2 => n20824, ZN => n25343);
   U18652 : OAI222_X1 port map( A1 => n20413, A2 => n23265, B1 => n20541, B2 =>
                           n23257, C1 => n20477, C2 => n23249, ZN => n25341);
   U18653 : NOR4_X1 port map( A1 => n25341, A2 => n16863, A3 => n16850, A4 => 
                           n16851, ZN => n25342);
   U18654 : AND3_X1 port map( A1 => n25344, A2 => n25343, A3 => n25342, ZN => 
                           n25345);
   U18655 : OAI222_X1 port map( A1 => n19517, A2 => n22936, B1 => n25345, B2 =>
                           n22799, C1 => n19645, C2 => n22516, ZN => n25346);
   U18656 : AOI221_X1 port map( B1 => n22922, B2 => n22140, C1 => n22971, C2 =>
                           n21148, A => n25346, ZN => n25354);
   U18657 : OAI22_X1 port map( A1 => n19133, A2 => n22976, B1 => n19261, B2 => 
                           n22633, ZN => n25347);
   U18658 : OAI222_X1 port map( A1 => n18941, A2 => n22952, B1 => n19197, B2 =>
                           n22966, C1 => n19069, C2 => n22637, ZN => n25348);
   U18659 : AOI221_X1 port map( B1 => n25391, B2 => n22182, C1 => n22962, C2 =>
                           n21264, A => n25348, ZN => n25352);
   U18660 : OAI22_X1 port map( A1 => n25394, A2 => n25349, B1 => n18685, B2 => 
                           n22947, ZN => n25350);
   U18661 : AOI221_X1 port map( B1 => n23280, B2 => n20953, C1 => n22494, C2 =>
                           n21693, A => n25350, ZN => n25351);
   U18662 : NAND4_X1 port map( A1 => n25352, A2 => n25353, A3 => n25351, A4 => 
                           n25354, ZN => n3336);
   U18663 : NAND2_X1 port map( A1 => n16827, A2 => n16828, ZN => n25356);
   U18664 : AOI21_X1 port map( B1 => n16831, B2 => n16832, A => n23201, ZN => 
                           n25355);
   U18665 : AOI221_X1 port map( B1 => n23217, B2 => n21876, C1 => n23209, C2 =>
                           n25356, A => n25355, ZN => n25360);
   U18666 : AOI222_X1 port map( A1 => n23241, A2 => n21319, B1 => n23233, B2 =>
                           n20995, C1 => n23225, C2 => n20802, ZN => n25359);
   U18667 : OAI222_X1 port map( A1 => n20475, A2 => n23265, B1 => n20603, B2 =>
                           n23257, C1 => n20539, C2 => n23249, ZN => n25357);
   U18668 : NOR4_X1 port map( A1 => n25357, A2 => n16836, A3 => n16823, A4 => 
                           n16824, ZN => n25358);
   U18669 : AND3_X1 port map( A1 => n25360, A2 => n25359, A3 => n25358, ZN => 
                           n25361);
   U18670 : OAI222_X1 port map( A1 => n19579, A2 => n22934, B1 => n25361, B2 =>
                           n22800, C1 => n19707, C2 => n22519, ZN => n25362);
   U18671 : AOI221_X1 port map( B1 => n22921, B2 => n22141, C1 => n22972, C2 =>
                           n21146, A => n25362, ZN => n25370);
   U18672 : OAI22_X1 port map( A1 => n19195, A2 => n22980, B1 => n19323, B2 => 
                           n22629, ZN => n25363);
   U18673 : AOI221_X1 port map( B1 => n22913, B2 => n22085, C1 => n22805, C2 =>
                           n21203, A => n25363, ZN => n25369);
   U18674 : OAI222_X1 port map( A1 => n19003, A2 => n22951, B1 => n19259, B2 =>
                           n22967, C1 => n19131, C2 => n22638, ZN => n25364);
   U18675 : AOI221_X1 port map( B1 => n25391, B2 => n22183, C1 => n22956, C2 =>
                           n21242, A => n25364, ZN => n25368);
   U18676 : OAI22_X1 port map( A1 => n25394, A2 => n25365, B1 => n18747, B2 => 
                           n22943, ZN => n25366);
   U18677 : AOI221_X1 port map( B1 => n23280, B2 => n20931, C1 => n22494, C2 =>
                           n21671, A => n25366, ZN => n25367);
   U18678 : NAND4_X1 port map( A1 => n25368, A2 => n25369, A3 => n25367, A4 => 
                           n25370, ZN => n3337);
   U18679 : NAND2_X1 port map( A1 => n16774, A2 => n16775, ZN => n25373);
   U18680 : AOI21_X1 port map( B1 => n16787, B2 => n16788, A => n23201, ZN => 
                           n25372);
   U18681 : AOI221_X1 port map( B1 => n23217, B2 => n21899, C1 => n23209, C2 =>
                           n25373, A => n25372, ZN => n25377);
   U18682 : AOI222_X1 port map( A1 => n23241, A2 => n21342, B1 => n23233, B2 =>
                           n21018, C1 => n23225, C2 => n20825, ZN => n25376);
   U18683 : OAI222_X1 port map( A1 => n20412, A2 => n23265, B1 => n20540, B2 =>
                           n23257, C1 => n20476, C2 => n23249, ZN => n25374);
   U18684 : NOR4_X1 port map( A1 => n25374, A2 => n16802, A3 => n16770, A4 => 
                           n16771, ZN => n25375);
   U18685 : AND3_X1 port map( A1 => n25377, A2 => n25376, A3 => n25375, ZN => 
                           n25380);
   U18686 : OAI222_X1 port map( A1 => n19516, A2 => n22934, B1 => n25380, B2 =>
                           n22799, C1 => n19644, C2 => n22520, ZN => n25382);
   U18687 : AOI221_X1 port map( B1 => n22922, B2 => n22142, C1 => n22973, C2 =>
                           n21149, A => n25382, ZN => n25399);
   U18688 : OAI22_X1 port map( A1 => n19132, A2 => n22979, B1 => n19260, B2 => 
                           n22642, ZN => n25386);
   U18689 : OAI222_X1 port map( A1 => n18940, A2 => n22955, B1 => n19196, B2 =>
                           n22967, C1 => n19068, C2 => n22639, ZN => n25390);
   U18690 : AOI221_X1 port map( B1 => n22801, B2 => n22057, C1 => n22962, C2 =>
                           n21265, A => n25390, ZN => n25397);
   U18691 : OAI22_X1 port map( A1 => n23270, A2 => n25393, B1 => n18684, B2 => 
                           n22944, ZN => n25395);
   U18692 : AOI221_X1 port map( B1 => n23280, B2 => n20954, C1 => n22494, C2 =>
                           n21694, A => n25395, ZN => n25396);
   U18693 : NAND4_X1 port map( A1 => n25396, A2 => n25398, A3 => n25397, A4 => 
                           n25399, ZN => n3338);

end SYN_BEHAVIORAL;
