
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_REGISTER_FILE is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_REGISTER_FILE;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_REGISTER_FILE.all;

entity REGISTER_FILE is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end REGISTER_FILE;

architecture SYN_BEHAVIORAL of REGISTER_FILE is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
      n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
      n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
      n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
      n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
      n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, 
      n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
      n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, 
      n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
      n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
      n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
      n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
      n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, 
      n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
      n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, 
      n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
      n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, 
      n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, 
      n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, 
      n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, 
      n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
      n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, 
      n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, 
      n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, 
      n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n4648, 
      n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, 
      n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, 
      n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, 
      n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, 
      n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, 
      n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, 
      n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, 
      n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, 
      n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, 
      n4739, n4740, n4741, n4742, n4743, n6741, n6742, n6743, n6744, n6745, 
      n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, 
      n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
      n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, 
      n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
      n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
      n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
      n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, 
      n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, 
      n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
      n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
      n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
      n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, 
      n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
      n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
      n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, 
      n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
      n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
      n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
      n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, 
      n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
      n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
      n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
      n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
      n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, 
      n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, 
      n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, 
      n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
      n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, 
      n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, 
      n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, 
      n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, 
      n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, 
      n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, 
      n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, 
      n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, 
      n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
      n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, 
      n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
      n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, 
      n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, 
      n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, 
      n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, 
      n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, 
      n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, 
      n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, 
      n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, 
      n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, 
      n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, 
      n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, 
      n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, 
      n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, 
      n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, 
      n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, 
      n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, 
      n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, 
      n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, 
      n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, 
      n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, 
      n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, 
      n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, 
      n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, 
      n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, 
      n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, 
      n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, 
      n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, 
      n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, 
      n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, 
      n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, 
      n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, 
      n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, 
      n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, 
      n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, 
      n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, 
      n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, 
      n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, 
      n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, 
      n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, 
      n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, 
      n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, 
      n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, 
      n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, 
      n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, 
      n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, 
      n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, 
      n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, 
      n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, 
      n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7654, n7655, n7656, 
      n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, 
      n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, 
      n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, 
      n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, 
      n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, 
      n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, 
      n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, 
      n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, 
      n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, 
      n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, 
      n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, 
      n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, 
      n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, 
      n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, 
      n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, 
      n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, 
      n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, 
      n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, 
      n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, 
      n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, 
      n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, 
      n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, 
      n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, 
      n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, 
      n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, 
      n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, 
      n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, 
      n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, 
      n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, 
      n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, 
      n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, 
      n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, 
      n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, 
      n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, 
      n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, 
      n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, 
      n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, 
      n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, 
      n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, 
      n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, 
      n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, 
      n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, 
      n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, 
      n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, 
      n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, 
      n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, 
      n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, 
      n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, 
      n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, 
      n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, 
      n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, 
      n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, 
      n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, 
      n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, 
      n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, 
      n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, 
      n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, 
      n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, 
      n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, 
      n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, 
      n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, 
      n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, 
      n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, 
      n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, 
      n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, 
      n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, 
      n8317, n8318, n8319, n8320, n8322, n8323, n8324, n8325, n8326, n8327, 
      n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, 
      n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, 
      n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, 
      n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, 
      n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, 
      n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, 
      n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, 
      n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, 
      n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, 
      n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, 
      n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, 
      n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, 
      n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, 
      n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, 
      n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, 
      n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, 
      n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, 
      n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, 
      n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
      n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, 
      n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, 
      n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, 
      n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, 
      n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, 
      n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, 
      n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, 
      n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, 
      n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, 
      n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, 
      n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, 
      n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, 
      n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, 
      n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, 
      n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, 
      n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, 
      n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, 
      n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, 
      n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, 
      n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, 
      n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, 
      n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, 
      n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, 
      n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, 
      n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, 
      n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, 
      n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, 
      n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, 
      n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, 
      n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, 
      n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, 
      n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, 
      n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, 
      n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, 
      n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, 
      n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, 
      n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, 
      n8888, n8889, n8890, n8891, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9084, n9085, n9086, n9087, 
      n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, 
      n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, 
      n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9148, n9149, 
      n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, 
      n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, 
      n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, 
      n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, 
      n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, 
      n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, 
      n9210, n9211, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, 
      n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, 
      n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, 
      n9272, n9273, n9274, n9275, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, 
      n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
      n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9404, n9405, 
      n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, 
      n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, 
      n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, 
      n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, 
      n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, 
      n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, 
      n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, 
      n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, 
      n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, 
      n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, 
      n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, 
      n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, 
      n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, 
      n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, 
      n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, 
      n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, 
      n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, 
      n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, 
      n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, 
      n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, 
      n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, 
      n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, 
      n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, 
      n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, 
      n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, 
      n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, 
      n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, 
      n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, 
      n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, 
      n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, 
      n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, 
      n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, 
      n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, 
      n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, 
      n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, 
      n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, 
      n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, 
      n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, 
      n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, 
      n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, 
      n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, 
      n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, 
      n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, 
      n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, 
      n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
      n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, 
      n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, 
      n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, 
      n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
      n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, 
      n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, 
      n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, 
      n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, 
      n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, 
      n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, 
      n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
      n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, 
      n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, 
      n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
      n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, 
      n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, 
      n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, 
      n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, 
      n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, 
      n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, 
      n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, 
      n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, 
      n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, 
      n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, 
      n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, 
      n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, 
      n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
      n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, 
      n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, 
      n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, 
      n10227, n10228, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639 : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT2_reg_31_inst : DFF_X1 port map( D => n2367, CK => CLK, Q => OUT2_31_port
                           , QN => n_1000);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2366, CK => CLK, Q => OUT2_30_port
                           , QN => n_1001);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2365, CK => CLK, Q => OUT2_29_port
                           , QN => n_1002);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2364, CK => CLK, Q => OUT2_28_port
                           , QN => n_1003);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2363, CK => CLK, Q => OUT2_27_port
                           , QN => n_1004);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2362, CK => CLK, Q => OUT2_26_port
                           , QN => n_1005);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2361, CK => CLK, Q => OUT2_25_port
                           , QN => n_1006);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2360, CK => CLK, Q => OUT2_24_port
                           , QN => n_1007);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2359, CK => CLK, Q => OUT2_23_port
                           , QN => n_1008);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2358, CK => CLK, Q => OUT2_22_port
                           , QN => n_1009);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2357, CK => CLK, Q => OUT2_21_port
                           , QN => n_1010);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2356, CK => CLK, Q => OUT2_20_port
                           , QN => n_1011);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2355, CK => CLK, Q => OUT2_19_port
                           , QN => n_1012);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2354, CK => CLK, Q => OUT2_18_port
                           , QN => n_1013);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2353, CK => CLK, Q => OUT2_17_port
                           , QN => n_1014);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2352, CK => CLK, Q => OUT2_16_port
                           , QN => n_1015);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2351, CK => CLK, Q => OUT2_15_port
                           , QN => n_1016);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2350, CK => CLK, Q => OUT2_14_port
                           , QN => n_1017);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2349, CK => CLK, Q => OUT2_13_port
                           , QN => n_1018);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2348, CK => CLK, Q => OUT2_12_port
                           , QN => n_1019);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2347, CK => CLK, Q => OUT2_11_port
                           , QN => n_1020);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2346, CK => CLK, Q => OUT2_10_port
                           , QN => n_1021);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2345, CK => CLK, Q => OUT2_9_port, 
                           QN => n_1022);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2344, CK => CLK, Q => OUT2_8_port, 
                           QN => n_1023);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2343, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1024);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2342, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1025);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2341, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1026);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2340, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1027);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2339, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1028);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2338, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1029);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2337, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1030);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2336, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1031);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => OUT1_14_port
                           , QN => n_1032);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => OUT1_13_port
                           , QN => n_1033);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => OUT1_12_port
                           , QN => n_1034);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => OUT1_11_port
                           , QN => n_1035);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => OUT1_10_port
                           , QN => n_1036);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => OUT1_9_port, 
                           QN => n_1037);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => OUT1_8_port, 
                           QN => n_1038);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => OUT1_7_port, 
                           QN => n_1039);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => OUT1_6_port, 
                           QN => n_1040);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => OUT1_5_port, 
                           QN => n_1041);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => OUT1_4_port, 
                           QN => n_1042);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => OUT1_3_port, 
                           QN => n_1043);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => OUT1_2_port, 
                           QN => n_1044);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => OUT1_1_port, 
                           QN => n_1045);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1046);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           n_1047, QN => n479);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           n_1048, QN => n478);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           n_1049, QN => n477);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           n_1050, QN => n476);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           n_1051, QN => n475);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           n_1052, QN => n474);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           n_1053, QN => n473);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           n_1054, QN => n472);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           n_1055, QN => n511);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           n_1056, QN => n510);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           n_1057, QN => n509);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           n_1058, QN => n508);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           n_1059, QN => n507);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           n_1060, QN => n506);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           n_1061, QN => n505);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           n_1062, QN => n504);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           n_1063, QN => n671);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           n_1064, QN => n670);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           n_1065, QN => n669);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           n_1066, QN => n668);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           n_1067, QN => n667);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           n_1068, QN => n666);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           n_1069, QN => n665);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           n_1070, QN => n664);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           n_1071, QN => n735);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           n_1072, QN => n734);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           n_1073, QN => n733);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           n_1074, QN => n732);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           n_1075, QN => n731);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           n_1076, QN => n730);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           n_1077, QN => n729);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           n_1078, QN => n728);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           n_1079, QN => n471);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           n_1080, QN => n470);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n_1081, QN => n469);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           n_1082, QN => n468);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n_1083, QN => n467);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           n_1084, QN => n466);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n_1085, QN => n465);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           n_1086, QN => n464);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           n_1087, QN => n503);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           n_1088, QN => n502);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n_1089, QN => n501);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           n_1090, QN => n500);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n_1091, QN => n499);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           n_1092, QN => n498);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n_1093, QN => n497);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           n_1094, QN => n496);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n_1095, QN => n495);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           n_1096, QN => n494);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n_1097, QN => n493);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           n_1098, QN => n492);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n_1099, QN => n491);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           n_1100, QN => n490);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n_1101, QN => n489);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           n_1102, QN => n488);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n_1103, QN => n487);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           n_1104, QN => n486);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n_1105, QN => n485);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           n_1106, QN => n484);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n_1107, QN => n483);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           n_1108, QN => n482);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n_1109, QN => n481);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           n_1110, QN => n480);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           n_1111, QN => n518);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n_1112, QN => n517);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           n_1113, QN => n516);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n_1114, QN => n515);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           n_1115, QN => n514);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n_1116, QN => n513);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           n_1117, QN => n512);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           n_1118, QN => n567);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n_1119, QN => n566);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n_1120, QN => n565);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           n_1121, QN => n564);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           n_1122, QN => n563);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           n_1123, QN => n562);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           n_1124, QN => n561);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           n_1125, QN => n560);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           n_1126, QN => n559);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           n_1127, QN => n558);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           n_1128, QN => n557);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           n_1129, QN => n556);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           n_1130, QN => n555);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n_1131, QN => n554);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n_1132, QN => n553);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n_1133, QN => n552);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n_1134, QN => n551);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n_1135, QN => n550);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n_1136, QN => n549);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n_1137, QN => n548);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n_1138, QN => n547);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n_1139, QN => n546);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           n_1140, QN => n545);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           n_1141, QN => n544);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n_1142, QN => n663);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n_1143, QN => n662);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n_1144, QN => n661);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n_1145, QN => n660);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n_1146, QN => n659);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n_1147, QN => n658);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n_1148, QN => n657);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n_1149, QN => n656);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n_1150, QN => n655);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n_1151, QN => n654);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n_1152, QN => n653);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n_1153, QN => n652);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n_1154, QN => n651);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n_1155, QN => n650);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n_1156, QN => n649);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n_1157, QN => n648);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n_1158, QN => n647);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n_1159, QN => n646);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           n_1160, QN => n645);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           n_1161, QN => n644);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           n_1162, QN => n643);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           n_1163, QN => n642);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           n_1164, QN => n641);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           n_1165, QN => n640);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n_1166, QN => n727);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n_1167, QN => n726);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n_1168, QN => n725);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n_1169, QN => n724);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n_1170, QN => n723);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n_1171, QN => n722);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n_1172, QN => n721);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n_1173, QN => n720);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n_1174, QN => n719);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n_1175, QN => n718);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n_1176, QN => n717);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n_1177, QN => n716);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n_1178, QN => n715);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n_1179, QN => n714);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n_1180, QN => n713);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n_1181, QN => n712);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n_1182, QN => n711);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n_1183, QN => n710);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           n_1184, QN => n709);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           n_1185, QN => n708);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           n_1186, QN => n707);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           n_1187, QN => n706);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           n_1188, QN => n705);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           n_1189, QN => n704);
   U7330 : NAND3_X1 port map( A1 => n8200, A2 => n10081, A3 => n8201, ZN => 
                           n7642);
   U7331 : NAND3_X1 port map( A1 => n8200, A2 => n10081, A3 => n8202, ZN => 
                           n7641);
   U7332 : NAND3_X1 port map( A1 => n8200, A2 => n10081, A3 => n8206, ZN => 
                           n7647);
   U7333 : NAND3_X1 port map( A1 => n8200, A2 => n10081, A3 => n8207, ZN => 
                           n7646);
   U7334 : NAND3_X1 port map( A1 => n8203, A2 => n10081, A3 => n8208, ZN => 
                           n7652);
   U7335 : NAND3_X1 port map( A1 => n8202, A2 => n10081, A3 => n8208, ZN => 
                           n7651);
   U7336 : NAND3_X1 port map( A1 => n8206, A2 => n10081, A3 => n8208, ZN => 
                           n7658);
   U7337 : NAND3_X1 port map( A1 => n8204, A2 => n10081, A3 => n8208, ZN => 
                           n7657);
   U7338 : NAND3_X1 port map( A1 => n8868, A2 => n9687, A3 => n8869, ZN => 
                           n8310);
   U7339 : NAND3_X1 port map( A1 => n8868, A2 => n9687, A3 => n8870, ZN => 
                           n8309);
   U7340 : NAND3_X1 port map( A1 => n8868, A2 => n9687, A3 => n8874, ZN => 
                           n8315);
   U7341 : NAND3_X1 port map( A1 => n8868, A2 => n9687, A3 => n8875, ZN => 
                           n8314);
   U7342 : NAND3_X1 port map( A1 => n8871, A2 => n9687, A3 => n8876, ZN => 
                           n8320);
   U7343 : NAND3_X1 port map( A1 => n8870, A2 => n9687, A3 => n8876, ZN => 
                           n8319);
   U7344 : NAND3_X1 port map( A1 => n8874, A2 => n9687, A3 => n8876, ZN => 
                           n8326);
   U7345 : NAND3_X1 port map( A1 => n8872, A2 => n9687, A3 => n8876, ZN => 
                           n8325);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           n7513, QN => n607);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           n7514, QN => n606);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           n7515, QN => n605);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           n7516, QN => n604);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n7517, QN => n603);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n7518, QN => n602);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n7519, QN => n601);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n7520, QN => n600);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n7609, QN => n599);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n7610, QN => n598);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n7611, QN => n597);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n7612, QN => n596);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n7613, QN => n595);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n7614, QN => n594);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n7615, QN => n593);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n7616, QN => n592);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n7617, QN => n591);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n7618, QN => n590);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n7619, QN => n589);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n7620, QN => n588);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n7621, QN => n587);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n7622, QN => n586);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => n7623
                           , QN => n585);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => n7624
                           , QN => n584);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => n7625
                           , QN => n583);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => n7626
                           , QN => n582);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => n7627
                           , QN => n581);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => n7628
                           , QN => n580);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => n7629
                           , QN => n579);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => n7630
                           , QN => n578);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => n7631
                           , QN => n577);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => n7632
                           , QN => n576);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           n_1190, QN => n543);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           n_1191, QN => n542);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           n_1192, QN => n541);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           n_1193, QN => n540);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           n_1194, QN => n539);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           n_1195, QN => n538);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           n_1196, QN => n537);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           n_1197, QN => n536);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           n_1198, QN => n575);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           n_1199, QN => n574);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           n_1200, QN => n573);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           n_1201, QN => n572);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           n_1202, QN => n571);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           n_1203, QN => n570);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           n_1204, QN => n569);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           n_1205, QN => n568);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           n_1206, QN => n535);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n_1207, QN => n534);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n_1208, QN => n533);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n_1209, QN => n532);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n_1210, QN => n531);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n_1211, QN => n530);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n_1212, QN => n529);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n_1213, QN => n528);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n_1214, QN => n527);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n_1215, QN => n526);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n_1216, QN => n525);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n_1217, QN => n524);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n_1218, QN => n523);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           n_1219, QN => n522);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n_1220, QN => n521);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           n_1221, QN => n520);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n_1222, QN => n519);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           n_1223, QN => n7234);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           n_1224, QN => n7235);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           n_1225, QN => n7236);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           n_1226, QN => n7237);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           n_1227, QN => n7238);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           n_1228, QN => n7239);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           n_1229, QN => n7240);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           n_1230, QN => n7241);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           n_1231, QN => n7010);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           n_1232, QN => n7011);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           n_1233, QN => n7012);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           n_1234, QN => n7013);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           n_1235, QN => n7014);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           n_1236, QN => n7015);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           n_1237, QN => n7016);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           n_1238, QN => n7017);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n_1239, QN => n7242);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n_1240, QN => n7243);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n_1241, QN => n7244);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           n_1242, QN => n7245);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           n_1243, QN => n7246);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           n_1244, QN => n7247);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           n_1245, QN => n7248);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           n_1246, QN => n7249);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           n_1247, QN => n7250);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           n_1248, QN => n7251);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           n_1249, QN => n7252);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           n_1250, QN => n7253);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           n_1251, QN => n7254);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n_1252, QN => n7255);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n_1253, QN => n7256);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n_1254, QN => n7257);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n_1255, QN => n7258);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n_1256, QN => n7259);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           n_1257, QN => n7260);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           n_1258, QN => n7261);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           n_1259, QN => n7262);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           n_1260, QN => n7263);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           n_1261, QN => n7264);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           n_1262, QN => n7265);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           n_1263, QN => n7018);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           n_1264, QN => n7019);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           n_1265, QN => n7020);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           n_1266, QN => n7021);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           n_1267, QN => n7022);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           n_1268, QN => n7023);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           n_1269, QN => n7024);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           n_1270, QN => n7025);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           n_1271, QN => n7026);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           n_1272, QN => n7027);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           n_1273, QN => n7028);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           n_1274, QN => n7029);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           n_1275, QN => n7030);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           n_1276, QN => n7031);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => n_1277
                           , QN => n7032);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => n_1278
                           , QN => n7033);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => n_1279
                           , QN => n7034);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => n_1280
                           , QN => n7035);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => n_1281
                           , QN => n7036);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => n_1282
                           , QN => n7037);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => n_1283
                           , QN => n7038);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => n_1284
                           , QN => n7039);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => n_1285
                           , QN => n7040);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => n_1286
                           , QN => n7041);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           n_1287, QN => n7393);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           n_1288, QN => n7394);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           n_1289, QN => n7395);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           n_1290, QN => n7396);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           n_1291, QN => n7397);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           n_1292, QN => n7398);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           n_1293, QN => n7399);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           n_1294, QN => n7400);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           n_1295, QN => n7361);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           n_1296, QN => n7362);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           n_1297, QN => n7363);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           n_1298, QN => n7364);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           n_1299, QN => n7365);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           n_1300, QN => n7366);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           n_1301, QN => n7367);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           n_1302, QN => n7368);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           n_1303, QN => n7329);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           n_1304, QN => n7330);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           n_1305, QN => n7331);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           n_1306, QN => n7332);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           n_1307, QN => n7333);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           n_1308, QN => n7334);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           n_1309, QN => n7335);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           n_1310, QN => n7336);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           n_1311, QN => n7074);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           n_1312, QN => n7075);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           n_1313, QN => n7076);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           n_1314, QN => n7077);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           n_1315, QN => n7078);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           n_1316, QN => n7079);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           n_1317, QN => n7080);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           n_1318, QN => n7081);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           n_1319, QN => n7202);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           n_1320, QN => n7203);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           n_1321, QN => n7204);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           n_1322, QN => n7205);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           n_1323, QN => n7206);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           n_1324, QN => n7207);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           n_1325, QN => n7208);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           n_1326, QN => n7209);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           n_1327, QN => n6978);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           n_1328, QN => n6979);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           n_1329, QN => n6980);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           n_1330, QN => n6981);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           n_1331, QN => n6982);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           n_1332, QN => n6983);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           n_1333, QN => n6984);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           n_1334, QN => n6985);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           n_1335, QN => n7425);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           n_1336, QN => n7426);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           n_1337, QN => n7427);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           n_1338, QN => n7428);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           n_1339, QN => n7429);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           n_1340, QN => n7430);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           n_1341, QN => n7431);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           n_1342, QN => n7432);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2335, CK => CLK, Q => 
                           n_1343, QN => n6786);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2334, CK => CLK, Q => 
                           n_1344, QN => n6787);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2333, CK => CLK, Q => 
                           n_1345, QN => n6788);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2332, CK => CLK, Q => 
                           n_1346, QN => n6789);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2331, CK => CLK, Q => 
                           n_1347, QN => n6790);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2330, CK => CLK, Q => 
                           n_1348, QN => n6791);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2329, CK => CLK, Q => 
                           n_1349, QN => n6792);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2328, CK => CLK, Q => 
                           n_1350, QN => n6793);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           n_1351, QN => n7401);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           n_1352, QN => n7402);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n_1353, QN => n7403);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           n_1354, QN => n7404);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n_1355, QN => n7405);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           n_1356, QN => n7406);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n_1357, QN => n7407);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           n_1358, QN => n7408);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n_1359, QN => n7409);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           n_1360, QN => n7410);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n_1361, QN => n7411);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           n_1362, QN => n7412);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n_1363, QN => n7413);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           n_1364, QN => n7414);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n_1365, QN => n7415);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           n_1366, QN => n7416);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n_1367, QN => n7417);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           n_1368, QN => n7418);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n_1369, QN => n7419);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           n_1370, QN => n7420);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n_1371, QN => n7421);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           n_1372, QN => n7422);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           n_1373, QN => n7423);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           n_1374, QN => n7424);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           n_1375, QN => n7369);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           n_1376, QN => n7370);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n_1377, QN => n7371);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           n_1378, QN => n7372);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n_1379, QN => n7373);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           n_1380, QN => n7374);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n_1381, QN => n7375);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           n_1382, QN => n7376);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n_1383, QN => n7377);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           n_1384, QN => n7378);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n_1385, QN => n7379);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           n_1386, QN => n7380);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n_1387, QN => n7381);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           n_1388, QN => n7382);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n_1389, QN => n7383);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           n_1390, QN => n7384);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n_1391, QN => n7385);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           n_1392, QN => n7386);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n_1393, QN => n7387);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           n_1394, QN => n7388);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n_1395, QN => n7389);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           n_1396, QN => n7390);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n_1397, QN => n7391);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           n_1398, QN => n7392);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           n_1399, QN => n7337);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n_1400, QN => n7338);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n_1401, QN => n7339);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n_1402, QN => n7340);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n_1403, QN => n7341);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n_1404, QN => n7342);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n_1405, QN => n7343);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n_1406, QN => n7344);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n_1407, QN => n7345);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n_1408, QN => n7346);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n_1409, QN => n7347);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n_1410, QN => n7348);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n_1411, QN => n7349);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n_1412, QN => n7350);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n_1413, QN => n7351);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n_1414, QN => n7352);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n_1415, QN => n7353);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n_1416, QN => n7354);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           n_1417, QN => n7355);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           n_1418, QN => n7356);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           n_1419, QN => n7357);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           n_1420, QN => n7358);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           n_1421, QN => n7359);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           n_1422, QN => n7360);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           n_1423, QN => n7082);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           n_1424, QN => n7083);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           n_1425, QN => n7084);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           n_1426, QN => n7085);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           n_1427, QN => n7086);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           n_1428, QN => n7087);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           n_1429, QN => n7088);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           n_1430, QN => n7089);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           n_1431, QN => n7090);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           n_1432, QN => n7091);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           n_1433, QN => n7092);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           n_1434, QN => n7093);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           n_1435, QN => n7094);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           n_1436, QN => n7095);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => n_1437
                           , QN => n7096);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => n_1438
                           , QN => n7097);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => n_1439
                           , QN => n7098);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => n_1440
                           , QN => n7099);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => n_1441
                           , QN => n7100);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => n_1442
                           , QN => n7101);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => n_1443
                           , QN => n7102);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => n_1444
                           , QN => n7103);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => n_1445
                           , QN => n7104);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => n_1446
                           , QN => n7105);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           n_1447, QN => n7106);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           n_1448, QN => n7107);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           n_1449, QN => n7108);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           n_1450, QN => n7109);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           n_1451, QN => n7110);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           n_1452, QN => n7111);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           n_1453, QN => n7112);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           n_1454, QN => n7113);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => 
                           n_1455, QN => n6946);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => 
                           n_1456, QN => n6947);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => 
                           n_1457, QN => n6948);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => 
                           n_1458, QN => n6949);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => 
                           n_1459, QN => n6950);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => 
                           n_1460, QN => n6951);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => 
                           n_1461, QN => n6952);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => 
                           n_1462, QN => n6953);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           n_1463, QN => n7210);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           n_1464, QN => n7211);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           n_1465, QN => n7212);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           n_1466, QN => n7213);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           n_1467, QN => n7214);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           n_1468, QN => n7215);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           n_1469, QN => n7216);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           n_1470, QN => n7217);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           n_1471, QN => n7218);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           n_1472, QN => n7219);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           n_1473, QN => n7220);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           n_1474, QN => n7221);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           n_1475, QN => n7222);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           n_1476, QN => n7223);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           n_1477, QN => n7224);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           n_1478, QN => n7225);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           n_1479, QN => n7226);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           n_1480, QN => n7227);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           n_1481, QN => n7228);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           n_1482, QN => n7229);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           n_1483, QN => n7230);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           n_1484, QN => n7231);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           n_1485, QN => n7232);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           n_1486, QN => n7233);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           n_1487, QN => n6986);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           n_1488, QN => n6987);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           n_1489, QN => n6988);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           n_1490, QN => n6989);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           n_1491, QN => n6990);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           n_1492, QN => n6991);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           n_1493, QN => n6992);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           n_1494, QN => n6993);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           n_1495, QN => n6994);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           n_1496, QN => n6995);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           n_1497, QN => n6996);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           n_1498, QN => n6997);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           n_1499, QN => n6998);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           n_1500, QN => n6999);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => n_1501
                           , QN => n7000);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => n_1502
                           , QN => n7001);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => n_1503
                           , QN => n7002);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => n_1504
                           , QN => n7003);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => n_1505
                           , QN => n7004);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => n_1506
                           , QN => n7005);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => n_1507
                           , QN => n7006);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => n_1508
                           , QN => n7007);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => n_1509
                           , QN => n7008);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => n_1510
                           , QN => n7009);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           n_1511, QN => n7433);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           n_1512, QN => n7434);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           n_1513, QN => n7435);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           n_1514, QN => n7436);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           n_1515, QN => n7437);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           n_1516, QN => n7438);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           n_1517, QN => n7439);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           n_1518, QN => n7440);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           n_1519, QN => n7441);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           n_1520, QN => n7442);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           n_1521, QN => n7443);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           n_1522, QN => n7444);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           n_1523, QN => n7445);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           n_1524, QN => n7446);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           n_1525, QN => n7447);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           n_1526, QN => n7448);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           n_1527, QN => n7449);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           n_1528, QN => n7450);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           n_1529, QN => n7451);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           n_1530, QN => n7452);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           n_1531, QN => n7453);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           n_1532, QN => n7454);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           n_1533, QN => n7455);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           n_1534, QN => n7456);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n_1535, QN => n7593);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           n_1536, QN => n7594);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n_1537, QN => n7595);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           n_1538, QN => n7596);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n_1539, QN => n7597);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           n_1540, QN => n7598);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n_1541, QN => n7599);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           n_1542, QN => n7600);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n_1543, QN => n7601);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           n_1544, QN => n7602);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n_1545, QN => n7603);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           n_1546, QN => n7604);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n_1547, QN => n7605);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           n_1548, QN => n7606);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           n_1549, QN => n7607);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           n_1550, QN => n7608);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2327, CK => CLK, Q => 
                           n_1551, QN => n6794);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2326, CK => CLK, Q => 
                           n_1552, QN => n6795);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2325, CK => CLK, Q => 
                           n_1553, QN => n6796);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2324, CK => CLK, Q => 
                           n_1554, QN => n6797);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2323, CK => CLK, Q => 
                           n_1555, QN => n6798);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2322, CK => CLK, Q => 
                           n_1556, QN => n6799);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2321, CK => CLK, Q => 
                           n_1557, QN => n6800);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2320, CK => CLK, Q => 
                           n_1558, QN => n6801);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2319, CK => CLK, Q => 
                           n_1559, QN => n6802);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2318, CK => CLK, Q => 
                           n_1560, QN => n6803);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2317, CK => CLK, Q => 
                           n_1561, QN => n6804);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2316, CK => CLK, Q => 
                           n_1562, QN => n6805);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2315, CK => CLK, Q => 
                           n_1563, QN => n6806);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2314, CK => CLK, Q => 
                           n_1564, QN => n6807);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2313, CK => CLK, Q => n_1565
                           , QN => n6808);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2312, CK => CLK, Q => n_1566
                           , QN => n6809);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2311, CK => CLK, Q => n_1567
                           , QN => n6810);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2310, CK => CLK, Q => n_1568
                           , QN => n6811);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2309, CK => CLK, Q => n_1569
                           , QN => n6812);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2308, CK => CLK, Q => n_1570
                           , QN => n6813);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2307, CK => CLK, Q => n_1571
                           , QN => n6814);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2306, CK => CLK, Q => n_1572
                           , QN => n6815);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2305, CK => CLK, Q => n_1573
                           , QN => n6816);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2304, CK => CLK, Q => n_1574
                           , QN => n6817);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           n_1575, QN => n7114);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           n_1576, QN => n7115);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           n_1577, QN => n7116);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           n_1578, QN => n7117);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           n_1579, QN => n7118);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           n_1580, QN => n7119);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           n_1581, QN => n7120);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           n_1582, QN => n7121);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           n_1583, QN => n7122);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           n_1584, QN => n7123);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           n_1585, QN => n7124);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           n_1586, QN => n7125);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           n_1587, QN => n7126);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           n_1588, QN => n7127);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           n_1589, QN => n7128);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           n_1590, QN => n7129);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           n_1591, QN => n7130);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           n_1592, QN => n7131);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           n_1593, QN => n7132);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           n_1594, QN => n7133);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           n_1595, QN => n7134);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           n_1596, QN => n7135);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           n_1597, QN => n7136);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           n_1598, QN => n7137);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => 
                           n_1599, QN => n6954);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           n_1600, QN => n6955);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           n_1601, QN => n6956);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           n_1602, QN => n6957);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           n_1603, QN => n6958);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           n_1604, QN => n6959);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           n_1605, QN => n6960);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           n_1606, QN => n6961);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           n_1607, QN => n6962);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           n_1608, QN => n6963);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           n_1609, QN => n6964);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           n_1610, QN => n6965);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           n_1611, QN => n6966);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           n_1612, QN => n6967);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => n_1613
                           , QN => n6968);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => n_1614
                           , QN => n6969);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => n_1615
                           , QN => n6970);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => n_1616
                           , QN => n6971);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => n_1617
                           , QN => n6972);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => n_1618
                           , QN => n6973);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => n_1619
                           , QN => n6974);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => n_1620
                           , QN => n6975);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => n_1621
                           , QN => n6976);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => n_1622
                           , QN => n6977);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           n4680, QN => n7497);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           n4681, QN => n7498);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           n4682, QN => n7499);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           n4683, QN => n7500);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           n4684, QN => n7501);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           n4685, QN => n7502);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           n4686, QN => n7503);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           n4687, QN => n7504);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n4648, QN => n7505);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           n4649, QN => n7506);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n4650, QN => n7507);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           n4651, QN => n7508);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n4652, QN => n7509);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           n4653, QN => n7510);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n4654, QN => n7511);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           n4655, QN => n7512);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           n9371, QN => n7633);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           n9370, QN => n7266);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           n9369, QN => n7267);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           n9368, QN => n7268);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n9367, QN => n7269);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n9366, QN => n7270);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n9365, QN => n7271);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n9364, QN => n7272);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => n9115
                           , QN => n7042);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => n9114
                           , QN => n7043);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => n9113
                           , QN => n7044);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => n9112
                           , QN => n7045);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => n9111
                           , QN => n7046);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => n9110
                           , QN => n7047);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => n9109
                           , QN => n7048);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => n9108
                           , QN => n7049);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2207, CK => CLK, Q => n9179
                           , QN => n6914);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2206, CK => CLK, Q => n9178
                           , QN => n6915);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2205, CK => CLK, Q => n9177
                           , QN => n6916);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2204, CK => CLK, Q => n9176
                           , QN => n6917);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => n9175
                           , QN => n6918);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => n9174
                           , QN => n6919);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => n9173
                           , QN => n6920);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => n9172
                           , QN => n6921);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2239, CK => CLK, Q => n9563
                           , QN => n6882);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2238, CK => CLK, Q => n9562
                           , QN => n6883);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2237, CK => CLK, Q => n9561
                           , QN => n6884);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2236, CK => CLK, Q => n9560
                           , QN => n6885);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2235, CK => CLK, Q => n9559
                           , QN => n6886);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2234, CK => CLK, Q => n9558
                           , QN => n6887);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2233, CK => CLK, Q => n9557
                           , QN => n6888);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2232, CK => CLK, Q => n9556
                           , QN => n6889);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           n4688, QN => n7545);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           n4689, QN => n7546);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           n4690, QN => n7547);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           n4691, QN => n7548);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           n4692, QN => n7549);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           n4693, QN => n7550);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           n4694, QN => n7551);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           n4695, QN => n7552);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           n4696, QN => n7553);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           n4697, QN => n7554);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           n4698, QN => n7555);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           n4699, QN => n7556);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           n4700, QN => n7557);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           n4701, QN => n7558);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n4702
                           , QN => n7559);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n4703
                           , QN => n7560);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n4704
                           , QN => n7561);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n4705
                           , QN => n7562);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n4706
                           , QN => n7563);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n4707
                           , QN => n7564);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n4708
                           , QN => n7565);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n4709
                           , QN => n7566);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n4710
                           , QN => n7567);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n4711
                           , QN => n7568);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n4656, QN => n7569);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           n4657, QN => n7570);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n4658, QN => n7571);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           n4659, QN => n7572);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n4660, QN => n7573);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           n4661, QN => n7574);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n4662, QN => n7575);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           n4663, QN => n7576);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n4664, QN => n7577);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           n4665, QN => n7578);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n4666, QN => n7579);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           n4667, QN => n7580);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n4668, QN => n7581);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           n4669, QN => n7582);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n4670
                           , QN => n7583);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n4671
                           , QN => n7584);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n4672
                           , QN => n7585);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n4673
                           , QN => n7586);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n4674
                           , QN => n7587);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n4675
                           , QN => n7588);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n4676
                           , QN => n7589);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n4677
                           , QN => n7590);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n4678
                           , QN => n7591);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n4679
                           , QN => n7592);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n9363, QN => n7273);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n9362, QN => n7274);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n9361, QN => n7275);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n9360, QN => n7276);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n9359, QN => n7277);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n9358, QN => n7278);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n9357, QN => n7279);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n9356, QN => n7280);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n9355, QN => n7281);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n9354, QN => n7282);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n9353, QN => n7283);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n9352, QN => n7284);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n9351, QN => n7285);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n9350, QN => n7286);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => n9349
                           , QN => n7287);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => n9348
                           , QN => n7288);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => n9347
                           , QN => n7289);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => n9346
                           , QN => n7290);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => n9345
                           , QN => n7291);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => n9344
                           , QN => n7292);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => n9343
                           , QN => n7293);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => n9342
                           , QN => n7294);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => n9341
                           , QN => n7295);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => n9340
                           , QN => n7296);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => n9107
                           , QN => n7050);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => n9106
                           , QN => n7051);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => n9105
                           , QN => n7052);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => n9104
                           , QN => n7053);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => n9103
                           , QN => n7054);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => n9102
                           , QN => n7055);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => n9101
                           , QN => n7056);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => n9100
                           , QN => n7057);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => n9099
                           , QN => n7058);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => n9098
                           , QN => n7059);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => n9097
                           , QN => n7060);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => n9096
                           , QN => n7061);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => n9095
                           , QN => n7062);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => n9094
                           , QN => n7063);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => n9093,
                           QN => n7064);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => n9092,
                           QN => n7065);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => n9091,
                           QN => n7066);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => n9090,
                           QN => n7067);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => n9089,
                           QN => n7068);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => n9088,
                           QN => n7069);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => n9087,
                           QN => n7070);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => n9086,
                           QN => n7071);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => n9085,
                           QN => n7072);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => n9084,
                           QN => n7073);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => n9171
                           , QN => n6922);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => n9170
                           , QN => n6923);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => n9169
                           , QN => n6924);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => n9168
                           , QN => n6925);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => n9167
                           , QN => n6926);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => n9166
                           , QN => n6927);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => n9165
                           , QN => n6928);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => n9164
                           , QN => n6929);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => n9163
                           , QN => n6930);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => n9162
                           , QN => n6931);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => n9161
                           , QN => n6932);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => n9160
                           , QN => n6933);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => n9159
                           , QN => n6934);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => n9158
                           , QN => n6935);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => n9157,
                           QN => n6936);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => n9156,
                           QN => n6937);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => n9155,
                           QN => n6938);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => n9154,
                           QN => n6939);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => n9153,
                           QN => n6940);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => n9152,
                           QN => n6941);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => n9151,
                           QN => n6942);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => n9150,
                           QN => n6943);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => n9149,
                           QN => n6944);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => n9148,
                           QN => n6945);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2231, CK => CLK, Q => n9555
                           , QN => n6890);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2230, CK => CLK, Q => n9554
                           , QN => n6891);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2229, CK => CLK, Q => n9553
                           , QN => n6892);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2228, CK => CLK, Q => n9552
                           , QN => n6893);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2227, CK => CLK, Q => n9551
                           , QN => n6894);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2226, CK => CLK, Q => n9550
                           , QN => n6895);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2225, CK => CLK, Q => n9549
                           , QN => n6896);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2224, CK => CLK, Q => n9548
                           , QN => n6897);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2223, CK => CLK, Q => n9547
                           , QN => n6898);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2222, CK => CLK, Q => n9546
                           , QN => n6899);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2221, CK => CLK, Q => n9545
                           , QN => n6900);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2220, CK => CLK, Q => n9544
                           , QN => n6901);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2219, CK => CLK, Q => n9543
                           , QN => n6902);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2218, CK => CLK, Q => n9542
                           , QN => n6903);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2217, CK => CLK, Q => n9541,
                           QN => n6904);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2216, CK => CLK, Q => n9540,
                           QN => n6905);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2215, CK => CLK, Q => n9539,
                           QN => n6906);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2214, CK => CLK, Q => n9538,
                           QN => n6907);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2213, CK => CLK, Q => n9537,
                           QN => n6908);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2212, CK => CLK, Q => n9536,
                           QN => n6909);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2211, CK => CLK, Q => n9535,
                           QN => n6910);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2210, CK => CLK, Q => n9534,
                           QN => n6911);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2209, CK => CLK, Q => n9533,
                           QN => n6912);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2208, CK => CLK, Q => n9532,
                           QN => n6913);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           n9275, QN => n7457);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           n9274, QN => n7458);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           n9273, QN => n7459);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           n9272, QN => n7460);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           n9271, QN => n7461);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           n9270, QN => n7462);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           n9269, QN => n7463);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           n9268, QN => n7464);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           n4712, QN => n7489);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           n4713, QN => n7490);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           n4714, QN => n7491);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           n4715, QN => n7492);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           n4716, QN => n7493);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           n4717, QN => n7494);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           n4718, QN => n7495);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           n4719, QN => n7496);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           n9339, QN => n7297);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           n9338, QN => n7298);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           n9337, QN => n7299);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           n9336, QN => n7300);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           n9335, QN => n7301);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           n9334, QN => n7302);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           n9333, QN => n7303);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           n9332, QN => n7304);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           n9051, QN => n7170);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           n9050, QN => n7171);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           n9049, QN => n7172);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           n9048, QN => n7173);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           n9047, QN => n7174);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           n9046, QN => n7175);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           n9045, QN => n7176);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           n9044, QN => n7177);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           n9435, QN => n7138);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           n9434, QN => n7139);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           n9433, QN => n7140);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           n9432, QN => n7141);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           n9431, QN => n7142);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           n9430, QN => n7143);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           n9429, QN => n7144);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           n9428, QN => n7145);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2271, CK => CLK, Q => n9595
                           , QN => n6850);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2270, CK => CLK, Q => n9594
                           , QN => n6851);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2269, CK => CLK, Q => n9593
                           , QN => n6852);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2268, CK => CLK, Q => n9592
                           , QN => n6853);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2267, CK => CLK, Q => n9591
                           , QN => n6854);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2266, CK => CLK, Q => n9590
                           , QN => n6855);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2265, CK => CLK, Q => n9589
                           , QN => n6856);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2264, CK => CLK, Q => n9588
                           , QN => n6857);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2303, CK => CLK, Q => n9211
                           , QN => n6818);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2302, CK => CLK, Q => n9210
                           , QN => n6819);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2301, CK => CLK, Q => n9209
                           , QN => n6820);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2300, CK => CLK, Q => n9208
                           , QN => n6821);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2299, CK => CLK, Q => n9207
                           , QN => n6822);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2298, CK => CLK, Q => n9206
                           , QN => n6823);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2297, CK => CLK, Q => n9205
                           , QN => n6824);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2296, CK => CLK, Q => n9204
                           , QN => n6825);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           n9267, QN => n7465);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           n9266, QN => n7466);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           n9265, QN => n7467);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           n9264, QN => n7468);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           n9263, QN => n7469);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           n9262, QN => n7470);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           n9261, QN => n7471);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           n9260, QN => n7472);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           n9259, QN => n7473);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           n9258, QN => n7474);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           n9257, QN => n7475);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           n9256, QN => n7476);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           n9255, QN => n7477);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           n9254, QN => n7478);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n9253
                           , QN => n7479);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n9252
                           , QN => n7480);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n9251
                           , QN => n7481);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n9250
                           , QN => n7482);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n9249
                           , QN => n7483);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n9248
                           , QN => n7484);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n9247
                           , QN => n7485);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n9246
                           , QN => n7486);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n9245
                           , QN => n7487);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n9244
                           , QN => n7488);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           n4720, QN => n7521);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           n4721, QN => n7522);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           n4722, QN => n7523);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           n4723, QN => n7524);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           n4724, QN => n7525);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           n4725, QN => n7526);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           n4726, QN => n7527);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           n4727, QN => n7528);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           n4728, QN => n7529);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           n4729, QN => n7530);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           n4730, QN => n7531);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           n4731, QN => n7532);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           n4732, QN => n7533);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           n4733, QN => n7534);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n4734
                           , QN => n7535);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n4735
                           , QN => n7536);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n4736
                           , QN => n7537);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n4737
                           , QN => n7538);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n4738
                           , QN => n7539);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n4739
                           , QN => n7540);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n4740
                           , QN => n7541);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n4741
                           , QN => n7542);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n4742
                           , QN => n7543);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n4743
                           , QN => n7544);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           n9331, QN => n7305);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n9330, QN => n7306);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n9329, QN => n7307);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n9328, QN => n7308);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n9327, QN => n7309);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n9326, QN => n7310);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n9325, QN => n7311);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n9324, QN => n7312);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n9323, QN => n7313);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n9322, QN => n7314);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n9321, QN => n7315);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n9320, QN => n7316);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n9319, QN => n7317);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n9318, QN => n7318);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => n9317
                           , QN => n7319);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => n9316
                           , QN => n7320);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => n9315
                           , QN => n7321);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => n9314
                           , QN => n7322);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => n9313
                           , QN => n7323);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => n9312
                           , QN => n7324);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => n9311
                           , QN => n7325);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => n9310
                           , QN => n7326);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => n9309
                           , QN => n7327);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => n9308
                           , QN => n7328);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n9043, QN => n7178);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n9042, QN => n7179);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n9041, QN => n7180);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           n9040, QN => n7181);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           n9039, QN => n7182);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           n9038, QN => n7183);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           n9037, QN => n7184);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           n9036, QN => n7185);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           n9035, QN => n7186);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           n9034, QN => n7187);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           n9033, QN => n7188);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           n9032, QN => n7189);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           n9031, QN => n7190);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           n9030, QN => n7191);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => n9029
                           , QN => n7192);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => n9028
                           , QN => n7193);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => n9027
                           , QN => n7194);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => n9026
                           , QN => n7195);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => n9025
                           , QN => n7196);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => n9024
                           , QN => n7197);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => n9023
                           , QN => n7198);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => n9022
                           , QN => n7199);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => n9021
                           , QN => n7200);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => n9020
                           , QN => n7201);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           n9427, QN => n7146);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           n9426, QN => n7147);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           n9425, QN => n7148);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           n9424, QN => n7149);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           n9423, QN => n7150);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           n9422, QN => n7151);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           n9421, QN => n7152);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           n9420, QN => n7153);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           n9419, QN => n7154);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           n9418, QN => n7155);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           n9417, QN => n7156);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           n9416, QN => n7157);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           n9415, QN => n7158);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           n9414, QN => n7159);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => n9413
                           , QN => n7160);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => n9412
                           , QN => n7161);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => n9411
                           , QN => n7162);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => n9410
                           , QN => n7163);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => n9409
                           , QN => n7164);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => n9408
                           , QN => n7165);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => n9407
                           , QN => n7166);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => n9406
                           , QN => n7167);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => n9405
                           , QN => n7168);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => n9404
                           , QN => n7169);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2263, CK => CLK, Q => n9587
                           , QN => n6858);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2262, CK => CLK, Q => n9586
                           , QN => n6859);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2261, CK => CLK, Q => n9585
                           , QN => n6860);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2260, CK => CLK, Q => n9584
                           , QN => n6861);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2259, CK => CLK, Q => n9583
                           , QN => n6862);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2258, CK => CLK, Q => n9582
                           , QN => n6863);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2257, CK => CLK, Q => n9581
                           , QN => n6864);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2256, CK => CLK, Q => n9580
                           , QN => n6865);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2255, CK => CLK, Q => n9579
                           , QN => n6866);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2254, CK => CLK, Q => n9578
                           , QN => n6867);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2253, CK => CLK, Q => n9577
                           , QN => n6868);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2252, CK => CLK, Q => n9576
                           , QN => n6869);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2251, CK => CLK, Q => n9575
                           , QN => n6870);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2250, CK => CLK, Q => n9574
                           , QN => n6871);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2249, CK => CLK, Q => n9573,
                           QN => n6872);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2248, CK => CLK, Q => n9572,
                           QN => n6873);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2247, CK => CLK, Q => n9571,
                           QN => n6874);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2246, CK => CLK, Q => n9570,
                           QN => n6875);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2245, CK => CLK, Q => n9569,
                           QN => n6876);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2244, CK => CLK, Q => n9568,
                           QN => n6877);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2243, CK => CLK, Q => n9567,
                           QN => n6878);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2242, CK => CLK, Q => n9566,
                           QN => n6879);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2241, CK => CLK, Q => n9565,
                           QN => n6880);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2240, CK => CLK, Q => n9564,
                           QN => n6881);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2295, CK => CLK, Q => n9203
                           , QN => n6826);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2294, CK => CLK, Q => n9202
                           , QN => n6827);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2293, CK => CLK, Q => n9201
                           , QN => n6828);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2292, CK => CLK, Q => n9200
                           , QN => n6829);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2291, CK => CLK, Q => n9199
                           , QN => n6830);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2290, CK => CLK, Q => n9198
                           , QN => n6831);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2289, CK => CLK, Q => n9197
                           , QN => n6832);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2288, CK => CLK, Q => n9196
                           , QN => n6833);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2287, CK => CLK, Q => n9195
                           , QN => n6834);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2286, CK => CLK, Q => n9194
                           , QN => n6835);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2285, CK => CLK, Q => n9193
                           , QN => n6836);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2284, CK => CLK, Q => n9192
                           , QN => n6837);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2283, CK => CLK, Q => n9191
                           , QN => n6838);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2282, CK => CLK, Q => n9190
                           , QN => n6839);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2281, CK => CLK, Q => n9189,
                           QN => n6840);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2280, CK => CLK, Q => n9188,
                           QN => n6841);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2279, CK => CLK, Q => n9187,
                           QN => n6842);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2278, CK => CLK, Q => n9186,
                           QN => n6843);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2277, CK => CLK, Q => n9185,
                           QN => n6844);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2276, CK => CLK, Q => n9184,
                           QN => n6845);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2275, CK => CLK, Q => n9183,
                           QN => n6846);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2274, CK => CLK, Q => n9182,
                           QN => n6847);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2273, CK => CLK, Q => n9181,
                           QN => n6848);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2272, CK => CLK, Q => n9180,
                           QN => n6849);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => OUT1_31_port
                           , QN => n_1623);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => OUT1_30_port
                           , QN => n_1624);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => OUT1_29_port
                           , QN => n_1625);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => OUT1_28_port
                           , QN => n_1626);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => OUT1_27_port
                           , QN => n_1627);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => OUT1_26_port
                           , QN => n_1628);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => OUT1_25_port
                           , QN => n_1629);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => OUT1_24_port
                           , QN => n_1630);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => OUT1_23_port
                           , QN => n_1631);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => OUT1_22_port
                           , QN => n_1632);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => OUT1_21_port
                           , QN => n_1633);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => OUT1_20_port
                           , QN => n_1634);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => OUT1_19_port
                           , QN => n_1635);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => OUT1_18_port
                           , QN => n_1636);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => OUT1_17_port
                           , QN => n_1637);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => OUT1_16_port
                           , QN => n_1638);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => OUT1_15_port
                           , QN => n_1639);
   U7346 : NOR2_X1 port map( A1 => n6745, A2 => ADD_WR(1), ZN => n8230);
   U7347 : NOR2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n8226);
   U7348 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n9596);
   U7349 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n9597);
   U7350 : BUF_X1 port map( A => n8266, Z => n9856);
   U7351 : BUF_X1 port map( A => n8271, Z => n9840);
   U7352 : BUF_X1 port map( A => n8276, Z => n9824);
   U7353 : BUF_X1 port map( A => n8279, Z => n9816);
   U7354 : BUF_X1 port map( A => n8281, Z => n9808);
   U7355 : BUF_X1 port map( A => n8283, Z => n9800);
   U7356 : BUF_X1 port map( A => n8285, Z => n9792);
   U7357 : BUF_X1 port map( A => n8290, Z => n9776);
   U7358 : BUF_X1 port map( A => n8297, Z => n9752);
   U7359 : BUF_X1 port map( A => n8299, Z => n9744);
   U7360 : BUF_X1 port map( A => n8301, Z => n9736);
   U7361 : BUF_X1 port map( A => n8294, Z => n9760);
   U7362 : BUF_X1 port map( A => n8292, Z => n9768);
   U7363 : BUF_X1 port map( A => n8288, Z => n9784);
   U7364 : BUF_X1 port map( A => n8273, Z => n9832);
   U7365 : BUF_X1 port map( A => n8269, Z => n9848);
   U7366 : BUF_X1 port map( A => n8264, Z => n9864);
   U7367 : BUF_X1 port map( A => n8262, Z => n9872);
   U7368 : BUF_X1 port map( A => n8260, Z => n9880);
   U7369 : BUF_X1 port map( A => n8257, Z => n9888);
   U7370 : BUF_X1 port map( A => n8255, Z => n9896);
   U7371 : BUF_X1 port map( A => n8253, Z => n9904);
   U7372 : BUF_X1 port map( A => n8251, Z => n9912);
   U7373 : BUF_X1 port map( A => n8248, Z => n9920);
   U7374 : BUF_X1 port map( A => n8246, Z => n9928);
   U7375 : BUF_X1 port map( A => n8244, Z => n9936);
   U7376 : BUF_X1 port map( A => n8242, Z => n9944);
   U7377 : BUF_X1 port map( A => n8239, Z => n9952);
   U7378 : BUF_X1 port map( A => n8235, Z => n9960);
   U7379 : BUF_X1 port map( A => n8232, Z => n9968);
   U7380 : BUF_X1 port map( A => n8229, Z => n9976);
   U7381 : BUF_X1 port map( A => n8225, Z => n9984);
   U7382 : BUF_X1 port map( A => n8319, Z => n9695);
   U7383 : BUF_X1 port map( A => n7651, Z => n10089);
   U7384 : BUF_X1 port map( A => n8320, Z => n9691);
   U7385 : BUF_X1 port map( A => n7652, Z => n10085);
   U7386 : BUF_X1 port map( A => n8326, Z => n9673);
   U7387 : BUF_X1 port map( A => n7658, Z => n10067);
   U7388 : BUF_X1 port map( A => n8325, Z => n9677);
   U7389 : BUF_X1 port map( A => n7657, Z => n10071);
   U7390 : BUF_X1 port map( A => n8314, Z => n9711);
   U7391 : BUF_X1 port map( A => n8315, Z => n9707);
   U7392 : BUF_X1 port map( A => n8309, Z => n9727);
   U7393 : BUF_X1 port map( A => n8310, Z => n9723);
   U7394 : BUF_X1 port map( A => n7646, Z => n10105);
   U7395 : BUF_X1 port map( A => n7647, Z => n10101);
   U7396 : BUF_X1 port map( A => n7641, Z => n10121);
   U7397 : BUF_X1 port map( A => n7642, Z => n10117);
   U7398 : BUF_X1 port map( A => n8311, Z => n9716);
   U7399 : BUF_X1 port map( A => n8312, Z => n9712);
   U7400 : BUF_X1 port map( A => n8316, Z => n9700);
   U7401 : BUF_X1 port map( A => n8317, Z => n9696);
   U7402 : BUF_X1 port map( A => n8306, Z => n9732);
   U7403 : BUF_X1 port map( A => n8307, Z => n9728);
   U7404 : BUF_X1 port map( A => n7644, Z => n10106);
   U7405 : BUF_X1 port map( A => n7643, Z => n10110);
   U7406 : BUF_X1 port map( A => n7649, Z => n10090);
   U7407 : BUF_X1 port map( A => n7648, Z => n10094);
   U7408 : BUF_X1 port map( A => n7639, Z => n10122);
   U7409 : BUF_X1 port map( A => n7638, Z => n10126);
   U7410 : BUF_X1 port map( A => n8351, Z => n9602);
   U7411 : BUF_X1 port map( A => n8352, Z => n9598);
   U7412 : BUF_X1 port map( A => n7683, Z => n9996);
   U7413 : BUF_X1 port map( A => n7684, Z => n9992);
   U7414 : BUF_X1 port map( A => n8331, Z => n9666);
   U7415 : BUF_X1 port map( A => n8332, Z => n9662);
   U7416 : BUF_X1 port map( A => n8342, Z => n9630);
   U7417 : BUF_X1 port map( A => n8343, Z => n9626);
   U7418 : BUF_X1 port map( A => n8337, Z => n9646);
   U7419 : BUF_X1 port map( A => n8338, Z => n9642);
   U7420 : BUF_X1 port map( A => n8348, Z => n9610);
   U7421 : BUF_X1 port map( A => n8349, Z => n9606);
   U7422 : BUF_X1 port map( A => n7664, Z => n10056);
   U7423 : BUF_X1 port map( A => n7663, Z => n10060);
   U7424 : BUF_X1 port map( A => n7675, Z => n10020);
   U7425 : BUF_X1 port map( A => n7674, Z => n10024);
   U7426 : BUF_X1 port map( A => n7670, Z => n10036);
   U7427 : BUF_X1 port map( A => n7669, Z => n10040);
   U7428 : BUF_X1 port map( A => n7681, Z => n10000);
   U7429 : BUF_X1 port map( A => n7680, Z => n10004);
   U7430 : BUF_X1 port map( A => n8270, Z => n9844);
   U7431 : BUF_X1 port map( A => n8280, Z => n9812);
   U7432 : BUF_X1 port map( A => n8282, Z => n9804);
   U7433 : BUF_X1 port map( A => n8289, Z => n9780);
   U7434 : BUF_X1 port map( A => n8298, Z => n9748);
   U7435 : BUF_X1 port map( A => n8300, Z => n9740);
   U7436 : BUF_X1 port map( A => n8291, Z => n9772);
   U7437 : BUF_X1 port map( A => n8272, Z => n9836);
   U7438 : BUF_X1 port map( A => n8263, Z => n9868);
   U7439 : BUF_X1 port map( A => n8261, Z => n9876);
   U7440 : BUF_X1 port map( A => n8254, Z => n9900);
   U7441 : BUF_X1 port map( A => n8252, Z => n9908);
   U7442 : BUF_X1 port map( A => n8245, Z => n9932);
   U7443 : BUF_X1 port map( A => n8243, Z => n9940);
   U7444 : BUF_X1 port map( A => n8234, Z => n9964);
   U7445 : BUF_X1 port map( A => n8231, Z => n9972);
   U7446 : BUF_X1 port map( A => n8336, Z => n9650);
   U7447 : BUF_X1 port map( A => n8335, Z => n9654);
   U7448 : BUF_X1 port map( A => n8334, Z => n9658);
   U7449 : BUF_X1 port map( A => n8347, Z => n9614);
   U7450 : BUF_X1 port map( A => n8346, Z => n9618);
   U7451 : BUF_X1 port map( A => n8345, Z => n9622);
   U7452 : BUF_X1 port map( A => n8340, Z => n9638);
   U7453 : BUF_X1 port map( A => n8341, Z => n9634);
   U7454 : BUF_X1 port map( A => n9596, Z => n9682);
   U7455 : BUF_X1 port map( A => n7668, Z => n10044);
   U7456 : BUF_X1 port map( A => n7667, Z => n10048);
   U7457 : BUF_X1 port map( A => n7666, Z => n10052);
   U7458 : BUF_X1 port map( A => n7679, Z => n10008);
   U7459 : BUF_X1 port map( A => n7678, Z => n10012);
   U7460 : BUF_X1 port map( A => n7677, Z => n10016);
   U7461 : BUF_X1 port map( A => n7673, Z => n10028);
   U7462 : BUF_X1 port map( A => n7672, Z => n10032);
   U7463 : BUF_X1 port map( A => n9597, Z => n10076);
   U7464 : BUF_X1 port map( A => n8265, Z => n9860);
   U7465 : BUF_X1 port map( A => n8275, Z => n9828);
   U7466 : BUF_X1 port map( A => n8278, Z => n9820);
   U7467 : BUF_X1 port map( A => n8284, Z => n9796);
   U7468 : BUF_X1 port map( A => n8296, Z => n9756);
   U7469 : BUF_X1 port map( A => n8293, Z => n9764);
   U7470 : BUF_X1 port map( A => n8287, Z => n9788);
   U7471 : BUF_X1 port map( A => n8268, Z => n9852);
   U7472 : BUF_X1 port map( A => n8259, Z => n9884);
   U7473 : BUF_X1 port map( A => n8256, Z => n9892);
   U7474 : BUF_X1 port map( A => n8250, Z => n9916);
   U7475 : BUF_X1 port map( A => n8247, Z => n9924);
   U7476 : BUF_X1 port map( A => n8241, Z => n9948);
   U7477 : BUF_X1 port map( A => n8238, Z => n9956);
   U7478 : BUF_X1 port map( A => n8228, Z => n9980);
   U7479 : BUF_X1 port map( A => n8224, Z => n9988);
   U7480 : BUF_X1 port map( A => n8323, Z => n9681);
   U7481 : BUF_X1 port map( A => n7655, Z => n10075);
   U7482 : BUF_X1 port map( A => n9856, Z => n9857);
   U7483 : BUF_X1 port map( A => n9856, Z => n9858);
   U7484 : BUF_X1 port map( A => n9840, Z => n9841);
   U7485 : BUF_X1 port map( A => n9840, Z => n9842);
   U7486 : BUF_X1 port map( A => n9824, Z => n9825);
   U7487 : BUF_X1 port map( A => n9824, Z => n9826);
   U7488 : BUF_X1 port map( A => n9816, Z => n9817);
   U7489 : BUF_X1 port map( A => n9816, Z => n9818);
   U7490 : BUF_X1 port map( A => n9808, Z => n9809);
   U7491 : BUF_X1 port map( A => n9808, Z => n9810);
   U7492 : BUF_X1 port map( A => n9800, Z => n9801);
   U7493 : BUF_X1 port map( A => n9800, Z => n9802);
   U7494 : BUF_X1 port map( A => n9792, Z => n9793);
   U7495 : BUF_X1 port map( A => n9792, Z => n9794);
   U7496 : BUF_X1 port map( A => n9776, Z => n9777);
   U7497 : BUF_X1 port map( A => n9776, Z => n9778);
   U7498 : BUF_X1 port map( A => n9752, Z => n9753);
   U7499 : BUF_X1 port map( A => n9752, Z => n9754);
   U7500 : BUF_X1 port map( A => n9744, Z => n9745);
   U7501 : BUF_X1 port map( A => n9744, Z => n9746);
   U7502 : BUF_X1 port map( A => n9736, Z => n9737);
   U7503 : BUF_X1 port map( A => n9736, Z => n9738);
   U7504 : BUF_X1 port map( A => n9760, Z => n9761);
   U7505 : BUF_X1 port map( A => n9760, Z => n9762);
   U7506 : BUF_X1 port map( A => n9768, Z => n9769);
   U7507 : BUF_X1 port map( A => n9768, Z => n9770);
   U7508 : BUF_X1 port map( A => n9784, Z => n9785);
   U7509 : BUF_X1 port map( A => n9784, Z => n9786);
   U7510 : BUF_X1 port map( A => n9832, Z => n9833);
   U7511 : BUF_X1 port map( A => n9832, Z => n9834);
   U7512 : BUF_X1 port map( A => n9848, Z => n9849);
   U7513 : BUF_X1 port map( A => n9848, Z => n9850);
   U7514 : BUF_X1 port map( A => n9864, Z => n9865);
   U7515 : BUF_X1 port map( A => n9864, Z => n9866);
   U7516 : BUF_X1 port map( A => n9872, Z => n9873);
   U7517 : BUF_X1 port map( A => n9872, Z => n9874);
   U7518 : BUF_X1 port map( A => n9880, Z => n9881);
   U7519 : BUF_X1 port map( A => n9880, Z => n9882);
   U7520 : BUF_X1 port map( A => n9888, Z => n9889);
   U7521 : BUF_X1 port map( A => n9888, Z => n9890);
   U7522 : BUF_X1 port map( A => n9896, Z => n9897);
   U7523 : BUF_X1 port map( A => n9896, Z => n9898);
   U7524 : BUF_X1 port map( A => n9904, Z => n9905);
   U7525 : BUF_X1 port map( A => n9904, Z => n9906);
   U7526 : BUF_X1 port map( A => n9912, Z => n9913);
   U7527 : BUF_X1 port map( A => n9912, Z => n9914);
   U7528 : BUF_X1 port map( A => n9920, Z => n9921);
   U7529 : BUF_X1 port map( A => n9920, Z => n9922);
   U7530 : BUF_X1 port map( A => n9928, Z => n9929);
   U7531 : BUF_X1 port map( A => n9928, Z => n9930);
   U7532 : BUF_X1 port map( A => n9936, Z => n9937);
   U7533 : BUF_X1 port map( A => n9936, Z => n9938);
   U7534 : BUF_X1 port map( A => n9944, Z => n9945);
   U7535 : BUF_X1 port map( A => n9944, Z => n9946);
   U7536 : BUF_X1 port map( A => n9952, Z => n9953);
   U7537 : BUF_X1 port map( A => n9952, Z => n9954);
   U7538 : BUF_X1 port map( A => n9960, Z => n9961);
   U7539 : BUF_X1 port map( A => n9960, Z => n9962);
   U7540 : BUF_X1 port map( A => n9968, Z => n9969);
   U7541 : BUF_X1 port map( A => n9968, Z => n9970);
   U7542 : BUF_X1 port map( A => n9976, Z => n9977);
   U7543 : BUF_X1 port map( A => n9976, Z => n9978);
   U7544 : BUF_X1 port map( A => n9984, Z => n9985);
   U7545 : BUF_X1 port map( A => n9984, Z => n9986);
   U7546 : BUF_X1 port map( A => n9856, Z => n9859);
   U7547 : BUF_X1 port map( A => n9840, Z => n9843);
   U7548 : BUF_X1 port map( A => n9824, Z => n9827);
   U7549 : BUF_X1 port map( A => n9816, Z => n9819);
   U7550 : BUF_X1 port map( A => n9808, Z => n9811);
   U7551 : BUF_X1 port map( A => n9800, Z => n9803);
   U7552 : BUF_X1 port map( A => n9792, Z => n9795);
   U7553 : BUF_X1 port map( A => n9776, Z => n9779);
   U7554 : BUF_X1 port map( A => n9752, Z => n9755);
   U7555 : BUF_X1 port map( A => n9744, Z => n9747);
   U7556 : BUF_X1 port map( A => n9736, Z => n9739);
   U7557 : BUF_X1 port map( A => n9760, Z => n9763);
   U7558 : BUF_X1 port map( A => n9768, Z => n9771);
   U7559 : BUF_X1 port map( A => n9784, Z => n9787);
   U7560 : BUF_X1 port map( A => n9832, Z => n9835);
   U7561 : BUF_X1 port map( A => n9848, Z => n9851);
   U7562 : BUF_X1 port map( A => n9864, Z => n9867);
   U7563 : BUF_X1 port map( A => n9872, Z => n9875);
   U7564 : BUF_X1 port map( A => n9880, Z => n9883);
   U7565 : BUF_X1 port map( A => n9888, Z => n9891);
   U7566 : BUF_X1 port map( A => n9896, Z => n9899);
   U7567 : BUF_X1 port map( A => n9904, Z => n9907);
   U7568 : BUF_X1 port map( A => n9912, Z => n9915);
   U7569 : BUF_X1 port map( A => n9920, Z => n9923);
   U7570 : BUF_X1 port map( A => n9928, Z => n9931);
   U7571 : BUF_X1 port map( A => n9936, Z => n9939);
   U7572 : BUF_X1 port map( A => n9944, Z => n9947);
   U7573 : BUF_X1 port map( A => n9952, Z => n9955);
   U7574 : BUF_X1 port map( A => n9960, Z => n9963);
   U7575 : BUF_X1 port map( A => n9968, Z => n9971);
   U7576 : BUF_X1 port map( A => n9976, Z => n9979);
   U7577 : BUF_X1 port map( A => n9984, Z => n9987);
   U7578 : NAND2_X1 port map( A1 => n10227, A2 => n9861, ZN => n8266);
   U7579 : NAND2_X1 port map( A1 => n10227, A2 => n9845, ZN => n8271);
   U7580 : NAND2_X1 port map( A1 => n10227, A2 => n9829, ZN => n8276);
   U7581 : NAND2_X1 port map( A1 => n10227, A2 => n9821, ZN => n8279);
   U7582 : NAND2_X1 port map( A1 => n10227, A2 => n9813, ZN => n8281);
   U7583 : NAND2_X1 port map( A1 => n10227, A2 => n9805, ZN => n8283);
   U7584 : NAND2_X1 port map( A1 => n10228, A2 => n9797, ZN => n8285);
   U7585 : NAND2_X1 port map( A1 => n10228, A2 => n9781, ZN => n8290);
   U7586 : NAND2_X1 port map( A1 => n10228, A2 => n9757, ZN => n8297);
   U7587 : NAND2_X1 port map( A1 => n10228, A2 => n9749, ZN => n8299);
   U7588 : NAND2_X1 port map( A1 => n10228, A2 => n9741, ZN => n8301);
   U7589 : NAND2_X1 port map( A1 => n10228, A2 => n9765, ZN => n8294);
   U7590 : NAND2_X1 port map( A1 => n10228, A2 => n9773, ZN => n8292);
   U7591 : NAND2_X1 port map( A1 => n10228, A2 => n9789, ZN => n8288);
   U7592 : NAND2_X1 port map( A1 => n10227, A2 => n9837, ZN => n8273);
   U7593 : NAND2_X1 port map( A1 => n10227, A2 => n9853, ZN => n8269);
   U7594 : NAND2_X1 port map( A1 => n10227, A2 => n9869, ZN => n8264);
   U7595 : NAND2_X1 port map( A1 => n10227, A2 => n9877, ZN => n8262);
   U7596 : NAND2_X1 port map( A1 => n10227, A2 => n9885, ZN => n8260);
   U7597 : NAND2_X1 port map( A1 => n10227, A2 => n9893, ZN => n8257);
   U7598 : NAND2_X1 port map( A1 => n10226, A2 => n9901, ZN => n8255);
   U7599 : NAND2_X1 port map( A1 => n10226, A2 => n9909, ZN => n8253);
   U7600 : NAND2_X1 port map( A1 => n10226, A2 => n9917, ZN => n8251);
   U7601 : NAND2_X1 port map( A1 => n10226, A2 => n9925, ZN => n8248);
   U7602 : NAND2_X1 port map( A1 => n10226, A2 => n9933, ZN => n8246);
   U7603 : NAND2_X1 port map( A1 => n10226, A2 => n9941, ZN => n8244);
   U7604 : NAND2_X1 port map( A1 => n10226, A2 => n9949, ZN => n8242);
   U7605 : NAND2_X1 port map( A1 => n10226, A2 => n9957, ZN => n8239);
   U7606 : NAND2_X1 port map( A1 => n10226, A2 => n9965, ZN => n8235);
   U7607 : NAND2_X1 port map( A1 => n10226, A2 => n9973, ZN => n8232);
   U7608 : NAND2_X1 port map( A1 => n10226, A2 => n9981, ZN => n8229);
   U7609 : NAND2_X1 port map( A1 => n10226, A2 => n9989, ZN => n8225);
   U7610 : BUF_X1 port map( A => n10089, Z => n10087);
   U7611 : BUF_X1 port map( A => n10056, Z => n10057);
   U7612 : BUF_X1 port map( A => n10020, Z => n10021);
   U7613 : BUF_X1 port map( A => n10036, Z => n10037);
   U7614 : BUF_X1 port map( A => n10000, Z => n10001);
   U7615 : BUF_X1 port map( A => n10056, Z => n10058);
   U7616 : BUF_X1 port map( A => n10020, Z => n10022);
   U7617 : BUF_X1 port map( A => n10036, Z => n10038);
   U7618 : BUF_X1 port map( A => n10000, Z => n10002);
   U7619 : BUF_X1 port map( A => n10106, Z => n10107);
   U7620 : BUF_X1 port map( A => n10090, Z => n10091);
   U7621 : BUF_X1 port map( A => n10122, Z => n10123);
   U7622 : BUF_X1 port map( A => n10106, Z => n10108);
   U7623 : BUF_X1 port map( A => n10090, Z => n10092);
   U7624 : BUF_X1 port map( A => n10122, Z => n10124);
   U7625 : BUF_X1 port map( A => n9988, Z => n9989);
   U7626 : BUF_X1 port map( A => n9988, Z => n9990);
   U7627 : BUF_X1 port map( A => n9677, Z => n9674);
   U7628 : BUF_X1 port map( A => n9711, Z => n9708);
   U7629 : BUF_X1 port map( A => n9695, Z => n9692);
   U7630 : BUF_X1 port map( A => n9727, Z => n9724);
   U7631 : BUF_X1 port map( A => n9677, Z => n9675);
   U7632 : BUF_X1 port map( A => n9711, Z => n9709);
   U7633 : BUF_X1 port map( A => n9695, Z => n9693);
   U7634 : BUF_X1 port map( A => n9727, Z => n9725);
   U7635 : BUF_X1 port map( A => n10105, Z => n10102);
   U7636 : BUF_X1 port map( A => n10121, Z => n10118);
   U7637 : BUF_X1 port map( A => n10105, Z => n10103);
   U7638 : BUF_X1 port map( A => n10121, Z => n10119);
   U7639 : BUF_X1 port map( A => n10089, Z => n10086);
   U7640 : BUF_X1 port map( A => n9860, Z => n9861);
   U7641 : BUF_X1 port map( A => n9844, Z => n9845);
   U7642 : BUF_X1 port map( A => n9828, Z => n9829);
   U7643 : BUF_X1 port map( A => n9820, Z => n9821);
   U7644 : BUF_X1 port map( A => n9812, Z => n9813);
   U7645 : BUF_X1 port map( A => n9804, Z => n9805);
   U7646 : BUF_X1 port map( A => n9796, Z => n9797);
   U7647 : BUF_X1 port map( A => n9780, Z => n9781);
   U7648 : BUF_X1 port map( A => n9756, Z => n9757);
   U7649 : BUF_X1 port map( A => n9748, Z => n9749);
   U7650 : BUF_X1 port map( A => n9740, Z => n9741);
   U7651 : BUF_X1 port map( A => n9764, Z => n9765);
   U7652 : BUF_X1 port map( A => n9772, Z => n9773);
   U7653 : BUF_X1 port map( A => n9788, Z => n9789);
   U7654 : BUF_X1 port map( A => n9836, Z => n9837);
   U7655 : BUF_X1 port map( A => n9852, Z => n9853);
   U7656 : BUF_X1 port map( A => n9868, Z => n9869);
   U7657 : BUF_X1 port map( A => n9876, Z => n9877);
   U7658 : BUF_X1 port map( A => n9884, Z => n9885);
   U7659 : BUF_X1 port map( A => n9892, Z => n9893);
   U7660 : BUF_X1 port map( A => n9900, Z => n9901);
   U7661 : BUF_X1 port map( A => n9908, Z => n9909);
   U7662 : BUF_X1 port map( A => n9916, Z => n9917);
   U7663 : BUF_X1 port map( A => n9924, Z => n9925);
   U7664 : BUF_X1 port map( A => n9932, Z => n9933);
   U7665 : BUF_X1 port map( A => n9940, Z => n9941);
   U7666 : BUF_X1 port map( A => n9948, Z => n9949);
   U7667 : BUF_X1 port map( A => n9956, Z => n9957);
   U7668 : BUF_X1 port map( A => n9964, Z => n9965);
   U7669 : BUF_X1 port map( A => n9972, Z => n9973);
   U7670 : BUF_X1 port map( A => n9980, Z => n9981);
   U7671 : BUF_X1 port map( A => n9638, Z => n9639);
   U7672 : BUF_X1 port map( A => n9602, Z => n9603);
   U7673 : BUF_X1 port map( A => n9638, Z => n9640);
   U7674 : BUF_X1 port map( A => n9602, Z => n9604);
   U7675 : BUF_X1 port map( A => n9996, Z => n9997);
   U7676 : BUF_X1 port map( A => n9996, Z => n9998);
   U7677 : BUF_X1 port map( A => n9860, Z => n9862);
   U7678 : BUF_X1 port map( A => n9844, Z => n9846);
   U7679 : BUF_X1 port map( A => n9828, Z => n9830);
   U7680 : BUF_X1 port map( A => n9820, Z => n9822);
   U7681 : BUF_X1 port map( A => n9812, Z => n9814);
   U7682 : BUF_X1 port map( A => n9804, Z => n9806);
   U7683 : BUF_X1 port map( A => n9796, Z => n9798);
   U7684 : BUF_X1 port map( A => n9780, Z => n9782);
   U7685 : BUF_X1 port map( A => n9756, Z => n9758);
   U7686 : BUF_X1 port map( A => n9748, Z => n9750);
   U7687 : BUF_X1 port map( A => n9740, Z => n9742);
   U7688 : BUF_X1 port map( A => n9764, Z => n9766);
   U7689 : BUF_X1 port map( A => n9772, Z => n9774);
   U7690 : BUF_X1 port map( A => n9788, Z => n9790);
   U7691 : BUF_X1 port map( A => n9836, Z => n9838);
   U7692 : BUF_X1 port map( A => n9852, Z => n9854);
   U7693 : BUF_X1 port map( A => n9868, Z => n9870);
   U7694 : BUF_X1 port map( A => n9876, Z => n9878);
   U7695 : BUF_X1 port map( A => n9884, Z => n9886);
   U7696 : BUF_X1 port map( A => n9892, Z => n9894);
   U7697 : BUF_X1 port map( A => n9900, Z => n9902);
   U7698 : BUF_X1 port map( A => n9908, Z => n9910);
   U7699 : BUF_X1 port map( A => n9916, Z => n9918);
   U7700 : BUF_X1 port map( A => n9924, Z => n9926);
   U7701 : BUF_X1 port map( A => n9932, Z => n9934);
   U7702 : BUF_X1 port map( A => n9940, Z => n9942);
   U7703 : BUF_X1 port map( A => n9948, Z => n9950);
   U7704 : BUF_X1 port map( A => n9956, Z => n9958);
   U7705 : BUF_X1 port map( A => n9964, Z => n9966);
   U7706 : BUF_X1 port map( A => n9972, Z => n9974);
   U7707 : BUF_X1 port map( A => n9980, Z => n9982);
   U7708 : BUF_X1 port map( A => n10044, Z => n10045);
   U7709 : BUF_X1 port map( A => n10008, Z => n10009);
   U7710 : BUF_X1 port map( A => n10044, Z => n10046);
   U7711 : BUF_X1 port map( A => n10008, Z => n10010);
   U7712 : BUF_X1 port map( A => n9673, Z => n9670);
   U7713 : BUF_X1 port map( A => n9707, Z => n9704);
   U7714 : BUF_X1 port map( A => n9691, Z => n9688);
   U7715 : BUF_X1 port map( A => n9723, Z => n9720);
   U7716 : BUF_X1 port map( A => n9673, Z => n9671);
   U7717 : BUF_X1 port map( A => n9707, Z => n9705);
   U7718 : BUF_X1 port map( A => n9691, Z => n9689);
   U7719 : BUF_X1 port map( A => n9723, Z => n9721);
   U7720 : BUF_X1 port map( A => n10117, Z => n10114);
   U7721 : BUF_X1 port map( A => n10117, Z => n10115);
   U7722 : BUF_X1 port map( A => n9634, Z => n9635);
   U7723 : BUF_X1 port map( A => n9598, Z => n9599);
   U7724 : BUF_X1 port map( A => n9634, Z => n9636);
   U7725 : BUF_X1 port map( A => n9598, Z => n9600);
   U7726 : BUF_X1 port map( A => n9992, Z => n9993);
   U7727 : BUF_X1 port map( A => n9992, Z => n9994);
   U7728 : BUF_X1 port map( A => n10048, Z => n10049);
   U7729 : BUF_X1 port map( A => n10012, Z => n10013);
   U7730 : BUF_X1 port map( A => n10048, Z => n10050);
   U7731 : BUF_X1 port map( A => n10012, Z => n10014);
   U7732 : BUF_X1 port map( A => n9682, Z => n9686);
   U7733 : BUF_X1 port map( A => n10076, Z => n10080);
   U7734 : BUF_X1 port map( A => n9682, Z => n9684);
   U7735 : BUF_X1 port map( A => n10076, Z => n10078);
   U7736 : BUF_X1 port map( A => n10052, Z => n10053);
   U7737 : BUF_X1 port map( A => n10016, Z => n10017);
   U7738 : BUF_X1 port map( A => n10052, Z => n10054);
   U7739 : BUF_X1 port map( A => n10016, Z => n10018);
   U7740 : BUF_X1 port map( A => n9666, Z => n9667);
   U7741 : BUF_X1 port map( A => n9630, Z => n9631);
   U7742 : BUF_X1 port map( A => n9646, Z => n9647);
   U7743 : BUF_X1 port map( A => n9610, Z => n9611);
   U7744 : BUF_X1 port map( A => n9666, Z => n9668);
   U7745 : BUF_X1 port map( A => n9630, Z => n9632);
   U7746 : BUF_X1 port map( A => n9646, Z => n9648);
   U7747 : BUF_X1 port map( A => n9610, Z => n9612);
   U7748 : BUF_X1 port map( A => n9716, Z => n9717);
   U7749 : BUF_X1 port map( A => n9700, Z => n9701);
   U7750 : BUF_X1 port map( A => n9732, Z => n9733);
   U7751 : BUF_X1 port map( A => n9716, Z => n9718);
   U7752 : BUF_X1 port map( A => n9700, Z => n9702);
   U7753 : BUF_X1 port map( A => n9732, Z => n9734);
   U7754 : BUF_X1 port map( A => n10126, Z => n10127);
   U7755 : BUF_X1 port map( A => n10126, Z => n10128);
   U7756 : BUF_X1 port map( A => n9682, Z => n9685);
   U7757 : BUF_X1 port map( A => n10076, Z => n10079);
   U7758 : BUF_X1 port map( A => n10067, Z => n10064);
   U7759 : BUF_X1 port map( A => n10101, Z => n10098);
   U7760 : BUF_X1 port map( A => n10085, Z => n10082);
   U7761 : BUF_X1 port map( A => n10067, Z => n10065);
   U7762 : BUF_X1 port map( A => n10101, Z => n10099);
   U7763 : BUF_X1 port map( A => n10085, Z => n10083);
   U7764 : BUF_X1 port map( A => n10028, Z => n10029);
   U7765 : BUF_X1 port map( A => n10028, Z => n10030);
   U7766 : BUF_X1 port map( A => n10071, Z => n10068);
   U7767 : BUF_X1 port map( A => n10071, Z => n10069);
   U7768 : BUF_X1 port map( A => n9662, Z => n9663);
   U7769 : BUF_X1 port map( A => n9626, Z => n9627);
   U7770 : BUF_X1 port map( A => n9642, Z => n9643);
   U7771 : BUF_X1 port map( A => n9606, Z => n9607);
   U7772 : BUF_X1 port map( A => n9662, Z => n9664);
   U7773 : BUF_X1 port map( A => n9626, Z => n9628);
   U7774 : BUF_X1 port map( A => n9642, Z => n9644);
   U7775 : BUF_X1 port map( A => n9606, Z => n9608);
   U7776 : BUF_X1 port map( A => n9712, Z => n9713);
   U7777 : BUF_X1 port map( A => n9696, Z => n9697);
   U7778 : BUF_X1 port map( A => n9728, Z => n9729);
   U7779 : BUF_X1 port map( A => n9712, Z => n9714);
   U7780 : BUF_X1 port map( A => n9696, Z => n9698);
   U7781 : BUF_X1 port map( A => n9728, Z => n9730);
   U7782 : BUF_X1 port map( A => n10060, Z => n10061);
   U7783 : BUF_X1 port map( A => n10024, Z => n10025);
   U7784 : BUF_X1 port map( A => n10040, Z => n10041);
   U7785 : BUF_X1 port map( A => n10004, Z => n10005);
   U7786 : BUF_X1 port map( A => n10060, Z => n10062);
   U7787 : BUF_X1 port map( A => n10024, Z => n10026);
   U7788 : BUF_X1 port map( A => n10040, Z => n10042);
   U7789 : BUF_X1 port map( A => n10004, Z => n10006);
   U7790 : BUF_X1 port map( A => n10110, Z => n10111);
   U7791 : BUF_X1 port map( A => n10094, Z => n10095);
   U7792 : BUF_X1 port map( A => n10110, Z => n10112);
   U7793 : BUF_X1 port map( A => n10094, Z => n10096);
   U7794 : BUF_X1 port map( A => n10032, Z => n10033);
   U7795 : BUF_X1 port map( A => n10032, Z => n10034);
   U7796 : BUF_X1 port map( A => n9650, Z => n9651);
   U7797 : BUF_X1 port map( A => n9614, Z => n9615);
   U7798 : BUF_X1 port map( A => n9650, Z => n9652);
   U7799 : BUF_X1 port map( A => n9614, Z => n9616);
   U7800 : BUF_X1 port map( A => n9654, Z => n9655);
   U7801 : BUF_X1 port map( A => n9618, Z => n9619);
   U7802 : BUF_X1 port map( A => n9654, Z => n9656);
   U7803 : BUF_X1 port map( A => n9618, Z => n9620);
   U7804 : BUF_X1 port map( A => n9658, Z => n9659);
   U7805 : BUF_X1 port map( A => n9622, Z => n9623);
   U7806 : BUF_X1 port map( A => n9658, Z => n9660);
   U7807 : BUF_X1 port map( A => n9622, Z => n9624);
   U7808 : BUF_X1 port map( A => n9860, Z => n9863);
   U7809 : BUF_X1 port map( A => n9844, Z => n9847);
   U7810 : BUF_X1 port map( A => n9828, Z => n9831);
   U7811 : BUF_X1 port map( A => n9820, Z => n9823);
   U7812 : BUF_X1 port map( A => n9812, Z => n9815);
   U7813 : BUF_X1 port map( A => n9804, Z => n9807);
   U7814 : BUF_X1 port map( A => n9796, Z => n9799);
   U7815 : BUF_X1 port map( A => n9780, Z => n9783);
   U7816 : BUF_X1 port map( A => n9756, Z => n9759);
   U7817 : BUF_X1 port map( A => n9748, Z => n9751);
   U7818 : BUF_X1 port map( A => n9740, Z => n9743);
   U7819 : BUF_X1 port map( A => n9764, Z => n9767);
   U7820 : BUF_X1 port map( A => n9772, Z => n9775);
   U7821 : BUF_X1 port map( A => n9788, Z => n9791);
   U7822 : BUF_X1 port map( A => n9836, Z => n9839);
   U7823 : BUF_X1 port map( A => n9852, Z => n9855);
   U7824 : BUF_X1 port map( A => n9868, Z => n9871);
   U7825 : BUF_X1 port map( A => n9876, Z => n9879);
   U7826 : BUF_X1 port map( A => n9884, Z => n9887);
   U7827 : BUF_X1 port map( A => n9892, Z => n9895);
   U7828 : BUF_X1 port map( A => n9900, Z => n9903);
   U7829 : BUF_X1 port map( A => n9908, Z => n9911);
   U7830 : BUF_X1 port map( A => n9916, Z => n9919);
   U7831 : BUF_X1 port map( A => n9924, Z => n9927);
   U7832 : BUF_X1 port map( A => n9932, Z => n9935);
   U7833 : BUF_X1 port map( A => n9940, Z => n9943);
   U7834 : BUF_X1 port map( A => n9948, Z => n9951);
   U7835 : BUF_X1 port map( A => n9956, Z => n9959);
   U7836 : BUF_X1 port map( A => n9964, Z => n9967);
   U7837 : BUF_X1 port map( A => n9972, Z => n9975);
   U7838 : BUF_X1 port map( A => n9980, Z => n9983);
   U7839 : BUF_X1 port map( A => n10056, Z => n10059);
   U7840 : BUF_X1 port map( A => n10020, Z => n10023);
   U7841 : BUF_X1 port map( A => n10036, Z => n10039);
   U7842 : BUF_X1 port map( A => n10000, Z => n10003);
   U7843 : BUF_X1 port map( A => n10106, Z => n10109);
   U7844 : BUF_X1 port map( A => n10090, Z => n10093);
   U7845 : BUF_X1 port map( A => n10122, Z => n10125);
   U7846 : BUF_X1 port map( A => n9677, Z => n9676);
   U7847 : BUF_X1 port map( A => n9711, Z => n9710);
   U7848 : BUF_X1 port map( A => n9695, Z => n9694);
   U7849 : BUF_X1 port map( A => n9727, Z => n9726);
   U7850 : BUF_X1 port map( A => n10105, Z => n10104);
   U7851 : BUF_X1 port map( A => n10121, Z => n10120);
   U7852 : BUF_X1 port map( A => n9638, Z => n9641);
   U7853 : BUF_X1 port map( A => n9602, Z => n9605);
   U7854 : BUF_X1 port map( A => n9996, Z => n9999);
   U7855 : BUF_X1 port map( A => n10044, Z => n10047);
   U7856 : BUF_X1 port map( A => n10008, Z => n10011);
   U7857 : BUF_X1 port map( A => n9673, Z => n9672);
   U7858 : BUF_X1 port map( A => n9707, Z => n9706);
   U7859 : BUF_X1 port map( A => n9691, Z => n9690);
   U7860 : BUF_X1 port map( A => n9723, Z => n9722);
   U7861 : BUF_X1 port map( A => n10117, Z => n10116);
   U7862 : BUF_X1 port map( A => n9634, Z => n9637);
   U7863 : BUF_X1 port map( A => n9598, Z => n9601);
   U7864 : BUF_X1 port map( A => n9992, Z => n9995);
   U7865 : BUF_X1 port map( A => n10048, Z => n10051);
   U7866 : BUF_X1 port map( A => n10012, Z => n10015);
   U7867 : BUF_X1 port map( A => n10052, Z => n10055);
   U7868 : BUF_X1 port map( A => n10016, Z => n10019);
   U7869 : BUF_X1 port map( A => n9666, Z => n9669);
   U7870 : BUF_X1 port map( A => n9630, Z => n9633);
   U7871 : BUF_X1 port map( A => n9646, Z => n9649);
   U7872 : BUF_X1 port map( A => n9610, Z => n9613);
   U7873 : BUF_X1 port map( A => n9716, Z => n9719);
   U7874 : BUF_X1 port map( A => n9700, Z => n9703);
   U7875 : BUF_X1 port map( A => n9732, Z => n9735);
   U7876 : BUF_X1 port map( A => n10126, Z => n10129);
   U7877 : BUF_X1 port map( A => n10067, Z => n10066);
   U7878 : BUF_X1 port map( A => n10101, Z => n10100);
   U7879 : BUF_X1 port map( A => n10085, Z => n10084);
   U7880 : BUF_X1 port map( A => n10071, Z => n10070);
   U7881 : BUF_X1 port map( A => n10028, Z => n10031);
   U7882 : BUF_X1 port map( A => n9662, Z => n9665);
   U7883 : BUF_X1 port map( A => n9626, Z => n9629);
   U7884 : BUF_X1 port map( A => n9642, Z => n9645);
   U7885 : BUF_X1 port map( A => n9606, Z => n9609);
   U7886 : BUF_X1 port map( A => n9712, Z => n9715);
   U7887 : BUF_X1 port map( A => n9696, Z => n9699);
   U7888 : BUF_X1 port map( A => n9728, Z => n9731);
   U7889 : BUF_X1 port map( A => n10060, Z => n10063);
   U7890 : BUF_X1 port map( A => n10024, Z => n10027);
   U7891 : BUF_X1 port map( A => n10040, Z => n10043);
   U7892 : BUF_X1 port map( A => n10004, Z => n10007);
   U7893 : BUF_X1 port map( A => n10110, Z => n10113);
   U7894 : BUF_X1 port map( A => n10094, Z => n10097);
   U7895 : BUF_X1 port map( A => n10032, Z => n10035);
   U7896 : BUF_X1 port map( A => n9650, Z => n9653);
   U7897 : BUF_X1 port map( A => n9614, Z => n9617);
   U7898 : BUF_X1 port map( A => n9654, Z => n9657);
   U7899 : BUF_X1 port map( A => n9618, Z => n9621);
   U7900 : BUF_X1 port map( A => n9658, Z => n9661);
   U7901 : BUF_X1 port map( A => n9622, Z => n9625);
   U7902 : BUF_X1 port map( A => n10089, Z => n10088);
   U7903 : BUF_X1 port map( A => n9988, Z => n9991);
   U7904 : OAI22_X1 port map( A1 => n10088, A2 => n7608, B1 => n10082, B2 => 
                           n7392, ZN => n8211);
   U7905 : OAI22_X1 port map( A1 => n10088, A2 => n7607, B1 => n10082, B2 => 
                           n7391, ZN => n8184);
   U7906 : OAI22_X1 port map( A1 => n10088, A2 => n7606, B1 => n10082, B2 => 
                           n7390, ZN => n8167);
   U7907 : OAI22_X1 port map( A1 => n10088, A2 => n7605, B1 => n10082, B2 => 
                           n7389, ZN => n8150);
   U7908 : OAI22_X1 port map( A1 => n10088, A2 => n7604, B1 => n10082, B2 => 
                           n7388, ZN => n8133);
   U7909 : OAI22_X1 port map( A1 => n10088, A2 => n7603, B1 => n10082, B2 => 
                           n7387, ZN => n8116);
   U7910 : OAI22_X1 port map( A1 => n10088, A2 => n7602, B1 => n10082, B2 => 
                           n7386, ZN => n8099);
   U7911 : OAI22_X1 port map( A1 => n10087, A2 => n7601, B1 => n10082, B2 => 
                           n7385, ZN => n8082);
   U7912 : OAI22_X1 port map( A1 => n10087, A2 => n7600, B1 => n10082, B2 => 
                           n7384, ZN => n8065);
   U7913 : OAI22_X1 port map( A1 => n10087, A2 => n7599, B1 => n10082, B2 => 
                           n7383, ZN => n8048);
   U7914 : OAI22_X1 port map( A1 => n10087, A2 => n7598, B1 => n10082, B2 => 
                           n7382, ZN => n8031);
   U7915 : OAI22_X1 port map( A1 => n10087, A2 => n7597, B1 => n10082, B2 => 
                           n7381, ZN => n8014);
   U7916 : OAI22_X1 port map( A1 => n10087, A2 => n7596, B1 => n10083, B2 => 
                           n7380, ZN => n7997);
   U7917 : OAI22_X1 port map( A1 => n10087, A2 => n7595, B1 => n10083, B2 => 
                           n7379, ZN => n7980);
   U7918 : OAI22_X1 port map( A1 => n10087, A2 => n7594, B1 => n10083, B2 => 
                           n7378, ZN => n7963);
   U7919 : OAI22_X1 port map( A1 => n10087, A2 => n7593, B1 => n10083, B2 => 
                           n7377, ZN => n7946);
   U7920 : OAI22_X1 port map( A1 => n7608, A2 => n9692, B1 => n7392, B2 => 
                           n9688, ZN => n8879);
   U7921 : OAI22_X1 port map( A1 => n7607, A2 => n9692, B1 => n7391, B2 => 
                           n9688, ZN => n8852);
   U7922 : OAI22_X1 port map( A1 => n7606, A2 => n9692, B1 => n7390, B2 => 
                           n9688, ZN => n8835);
   U7923 : OAI22_X1 port map( A1 => n7605, A2 => n9692, B1 => n7389, B2 => 
                           n9688, ZN => n8818);
   U7924 : OAI22_X1 port map( A1 => n7604, A2 => n9692, B1 => n7388, B2 => 
                           n9688, ZN => n8801);
   U7925 : OAI22_X1 port map( A1 => n7603, A2 => n9692, B1 => n7387, B2 => 
                           n9688, ZN => n8784);
   U7926 : OAI22_X1 port map( A1 => n7602, A2 => n9692, B1 => n7386, B2 => 
                           n9688, ZN => n8767);
   U7927 : OAI22_X1 port map( A1 => n7601, A2 => n9692, B1 => n7385, B2 => 
                           n9688, ZN => n8750);
   U7928 : OAI22_X1 port map( A1 => n7600, A2 => n9692, B1 => n7384, B2 => 
                           n9688, ZN => n8733);
   U7929 : OAI22_X1 port map( A1 => n7599, A2 => n9692, B1 => n7383, B2 => 
                           n9688, ZN => n8716);
   U7930 : OAI22_X1 port map( A1 => n7598, A2 => n9692, B1 => n7382, B2 => 
                           n9688, ZN => n8699);
   U7931 : OAI22_X1 port map( A1 => n7597, A2 => n9692, B1 => n7381, B2 => 
                           n9688, ZN => n8682);
   U7932 : OAI22_X1 port map( A1 => n7596, A2 => n9693, B1 => n7380, B2 => 
                           n9689, ZN => n8665);
   U7933 : OAI22_X1 port map( A1 => n7595, A2 => n9693, B1 => n7379, B2 => 
                           n9689, ZN => n8648);
   U7934 : OAI22_X1 port map( A1 => n7594, A2 => n9693, B1 => n7378, B2 => 
                           n9689, ZN => n8631);
   U7935 : OAI22_X1 port map( A1 => n7593, A2 => n9693, B1 => n7377, B2 => 
                           n9689, ZN => n8614);
   U7936 : OAI22_X1 port map( A1 => n10131, A2 => n9797, B1 => n7608, B2 => 
                           n9793, ZN => n1536);
   U7937 : OAI22_X1 port map( A1 => n10134, A2 => n9797, B1 => n7607, B2 => 
                           n9793, ZN => n1537);
   U7938 : OAI22_X1 port map( A1 => n10137, A2 => n9797, B1 => n7606, B2 => 
                           n9793, ZN => n1538);
   U7939 : OAI22_X1 port map( A1 => n10140, A2 => n9797, B1 => n7605, B2 => 
                           n9793, ZN => n1539);
   U7940 : OAI22_X1 port map( A1 => n10143, A2 => n9797, B1 => n7604, B2 => 
                           n9793, ZN => n1540);
   U7941 : OAI22_X1 port map( A1 => n10146, A2 => n9797, B1 => n7603, B2 => 
                           n9793, ZN => n1541);
   U7942 : OAI22_X1 port map( A1 => n10149, A2 => n9797, B1 => n7602, B2 => 
                           n9793, ZN => n1542);
   U7943 : OAI22_X1 port map( A1 => n10152, A2 => n9797, B1 => n7601, B2 => 
                           n9793, ZN => n1543);
   U7944 : OAI22_X1 port map( A1 => n10155, A2 => n9797, B1 => n7600, B2 => 
                           n9793, ZN => n1544);
   U7945 : OAI22_X1 port map( A1 => n10158, A2 => n9797, B1 => n7599, B2 => 
                           n9793, ZN => n1545);
   U7946 : OAI22_X1 port map( A1 => n10161, A2 => n9797, B1 => n7598, B2 => 
                           n9793, ZN => n1546);
   U7947 : OAI22_X1 port map( A1 => n10164, A2 => n9798, B1 => n7597, B2 => 
                           n9793, ZN => n1547);
   U7948 : OAI22_X1 port map( A1 => n10167, A2 => n9798, B1 => n7596, B2 => 
                           n9794, ZN => n1548);
   U7949 : OAI22_X1 port map( A1 => n10170, A2 => n9798, B1 => n7595, B2 => 
                           n9794, ZN => n1549);
   U7950 : OAI22_X1 port map( A1 => n10173, A2 => n9798, B1 => n7594, B2 => 
                           n9794, ZN => n1550);
   U7951 : OAI22_X1 port map( A1 => n10176, A2 => n9798, B1 => n7593, B2 => 
                           n9794, ZN => n1551);
   U7952 : OAI22_X1 port map( A1 => n10132, A2 => n9765, B1 => n7456, B2 => 
                           n9761, ZN => n1408);
   U7953 : OAI22_X1 port map( A1 => n10135, A2 => n9765, B1 => n7455, B2 => 
                           n9761, ZN => n1409);
   U7954 : OAI22_X1 port map( A1 => n10138, A2 => n9765, B1 => n7454, B2 => 
                           n9761, ZN => n1410);
   U7955 : OAI22_X1 port map( A1 => n10141, A2 => n9765, B1 => n7453, B2 => 
                           n9761, ZN => n1411);
   U7956 : OAI22_X1 port map( A1 => n10144, A2 => n9765, B1 => n7452, B2 => 
                           n9761, ZN => n1412);
   U7957 : OAI22_X1 port map( A1 => n10147, A2 => n9765, B1 => n7451, B2 => 
                           n9761, ZN => n1413);
   U7958 : OAI22_X1 port map( A1 => n10150, A2 => n9765, B1 => n7450, B2 => 
                           n9761, ZN => n1414);
   U7959 : OAI22_X1 port map( A1 => n10153, A2 => n9765, B1 => n7449, B2 => 
                           n9761, ZN => n1415);
   U7960 : OAI22_X1 port map( A1 => n10156, A2 => n9765, B1 => n7448, B2 => 
                           n9761, ZN => n1416);
   U7961 : OAI22_X1 port map( A1 => n10159, A2 => n9765, B1 => n7447, B2 => 
                           n9761, ZN => n1417);
   U7962 : OAI22_X1 port map( A1 => n10162, A2 => n9765, B1 => n7446, B2 => 
                           n9761, ZN => n1418);
   U7963 : OAI22_X1 port map( A1 => n10165, A2 => n9766, B1 => n7445, B2 => 
                           n9761, ZN => n1419);
   U7964 : OAI22_X1 port map( A1 => n10168, A2 => n9766, B1 => n7444, B2 => 
                           n9762, ZN => n1420);
   U7965 : OAI22_X1 port map( A1 => n10171, A2 => n9766, B1 => n7443, B2 => 
                           n9762, ZN => n1421);
   U7966 : OAI22_X1 port map( A1 => n10174, A2 => n9766, B1 => n7442, B2 => 
                           n9762, ZN => n1422);
   U7967 : OAI22_X1 port map( A1 => n10177, A2 => n9766, B1 => n7441, B2 => 
                           n9762, ZN => n1423);
   U7968 : OAI22_X1 port map( A1 => n10180, A2 => n9766, B1 => n7440, B2 => 
                           n9762, ZN => n1424);
   U7969 : OAI22_X1 port map( A1 => n10183, A2 => n9766, B1 => n7439, B2 => 
                           n9762, ZN => n1425);
   U7970 : OAI22_X1 port map( A1 => n10186, A2 => n9766, B1 => n7438, B2 => 
                           n9762, ZN => n1426);
   U7971 : OAI22_X1 port map( A1 => n10189, A2 => n9766, B1 => n7437, B2 => 
                           n9762, ZN => n1427);
   U7972 : OAI22_X1 port map( A1 => n10192, A2 => n9766, B1 => n7436, B2 => 
                           n9762, ZN => n1428);
   U7973 : OAI22_X1 port map( A1 => n10195, A2 => n9766, B1 => n7435, B2 => 
                           n9762, ZN => n1429);
   U7974 : OAI22_X1 port map( A1 => n10198, A2 => n9766, B1 => n7434, B2 => 
                           n9762, ZN => n1430);
   U7975 : OAI22_X1 port map( A1 => n10201, A2 => n9767, B1 => n7433, B2 => 
                           n9762, ZN => n1431);
   U7976 : OAI22_X1 port map( A1 => n10204, A2 => n9767, B1 => n7432, B2 => 
                           n9763, ZN => n1432);
   U7977 : OAI22_X1 port map( A1 => n10207, A2 => n9767, B1 => n7431, B2 => 
                           n9763, ZN => n1433);
   U7978 : OAI22_X1 port map( A1 => n10210, A2 => n9767, B1 => n7430, B2 => 
                           n9763, ZN => n1434);
   U7979 : OAI22_X1 port map( A1 => n10213, A2 => n9767, B1 => n7429, B2 => 
                           n9763, ZN => n1435);
   U7980 : OAI22_X1 port map( A1 => n10216, A2 => n9767, B1 => n7428, B2 => 
                           n9763, ZN => n1436);
   U7981 : OAI22_X1 port map( A1 => n10219, A2 => n9767, B1 => n7427, B2 => 
                           n9763, ZN => n1437);
   U7982 : OAI22_X1 port map( A1 => n10222, A2 => n9767, B1 => n7426, B2 => 
                           n9763, ZN => n1438);
   U7983 : OAI22_X1 port map( A1 => n10225, A2 => n9767, B1 => n7425, B2 => 
                           n9763, ZN => n1439);
   U7984 : OAI22_X1 port map( A1 => n9989, A2 => n10130, B1 => n6817, B2 => 
                           n9985, ZN => n2304);
   U7985 : OAI22_X1 port map( A1 => n9989, A2 => n10133, B1 => n6816, B2 => 
                           n9985, ZN => n2305);
   U7986 : OAI22_X1 port map( A1 => n9989, A2 => n10136, B1 => n6815, B2 => 
                           n9985, ZN => n2306);
   U7987 : OAI22_X1 port map( A1 => n9989, A2 => n10139, B1 => n6814, B2 => 
                           n9985, ZN => n2307);
   U7988 : OAI22_X1 port map( A1 => n9989, A2 => n10142, B1 => n6813, B2 => 
                           n9985, ZN => n2308);
   U7989 : OAI22_X1 port map( A1 => n9989, A2 => n10145, B1 => n6812, B2 => 
                           n9985, ZN => n2309);
   U7990 : OAI22_X1 port map( A1 => n9989, A2 => n10148, B1 => n6811, B2 => 
                           n9985, ZN => n2310);
   U7991 : OAI22_X1 port map( A1 => n9989, A2 => n10151, B1 => n6810, B2 => 
                           n9985, ZN => n2311);
   U7992 : OAI22_X1 port map( A1 => n9989, A2 => n10154, B1 => n6809, B2 => 
                           n9985, ZN => n2312);
   U7993 : OAI22_X1 port map( A1 => n9989, A2 => n10157, B1 => n6808, B2 => 
                           n9985, ZN => n2313);
   U7994 : OAI22_X1 port map( A1 => n9989, A2 => n10160, B1 => n6807, B2 => 
                           n9985, ZN => n2314);
   U7995 : OAI22_X1 port map( A1 => n9989, A2 => n10163, B1 => n6806, B2 => 
                           n9985, ZN => n2315);
   U7996 : OAI22_X1 port map( A1 => n9990, A2 => n10166, B1 => n6805, B2 => 
                           n9986, ZN => n2316);
   U7997 : OAI22_X1 port map( A1 => n9990, A2 => n10169, B1 => n6804, B2 => 
                           n9986, ZN => n2317);
   U7998 : OAI22_X1 port map( A1 => n9990, A2 => n10172, B1 => n6803, B2 => 
                           n9986, ZN => n2318);
   U7999 : OAI22_X1 port map( A1 => n9990, A2 => n10175, B1 => n6802, B2 => 
                           n9986, ZN => n2319);
   U8000 : OAI22_X1 port map( A1 => n9990, A2 => n10178, B1 => n6801, B2 => 
                           n9986, ZN => n2320);
   U8001 : OAI22_X1 port map( A1 => n9990, A2 => n10181, B1 => n6800, B2 => 
                           n9986, ZN => n2321);
   U8002 : OAI22_X1 port map( A1 => n9990, A2 => n10184, B1 => n6799, B2 => 
                           n9986, ZN => n2322);
   U8003 : OAI22_X1 port map( A1 => n9990, A2 => n10187, B1 => n6798, B2 => 
                           n9986, ZN => n2323);
   U8004 : OAI22_X1 port map( A1 => n9990, A2 => n10190, B1 => n6797, B2 => 
                           n9986, ZN => n2324);
   U8005 : OAI22_X1 port map( A1 => n9990, A2 => n10193, B1 => n6796, B2 => 
                           n9986, ZN => n2325);
   U8006 : OAI22_X1 port map( A1 => n9990, A2 => n10196, B1 => n6795, B2 => 
                           n9986, ZN => n2326);
   U8007 : OAI22_X1 port map( A1 => n9990, A2 => n10199, B1 => n6794, B2 => 
                           n9986, ZN => n2327);
   U8008 : OAI22_X1 port map( A1 => n9990, A2 => n10202, B1 => n6793, B2 => 
                           n9987, ZN => n2328);
   U8009 : OAI22_X1 port map( A1 => n9991, A2 => n10205, B1 => n6792, B2 => 
                           n9987, ZN => n2329);
   U8010 : OAI22_X1 port map( A1 => n9991, A2 => n10208, B1 => n6791, B2 => 
                           n9987, ZN => n2330);
   U8011 : OAI22_X1 port map( A1 => n9991, A2 => n10211, B1 => n6790, B2 => 
                           n9987, ZN => n2331);
   U8012 : OAI22_X1 port map( A1 => n9991, A2 => n10214, B1 => n6789, B2 => 
                           n9987, ZN => n2332);
   U8013 : OAI22_X1 port map( A1 => n9991, A2 => n10217, B1 => n6788, B2 => 
                           n9987, ZN => n2333);
   U8014 : OAI22_X1 port map( A1 => n9991, A2 => n10220, B1 => n6787, B2 => 
                           n9987, ZN => n2334);
   U8015 : OAI22_X1 port map( A1 => n9991, A2 => n10223, B1 => n6786, B2 => 
                           n9987, ZN => n2335);
   U8016 : OAI22_X1 port map( A1 => n10131, A2 => n9885, B1 => n7233, B2 => 
                           n9881, ZN => n1888);
   U8017 : OAI22_X1 port map( A1 => n10134, A2 => n9885, B1 => n7232, B2 => 
                           n9881, ZN => n1889);
   U8018 : OAI22_X1 port map( A1 => n10137, A2 => n9885, B1 => n7231, B2 => 
                           n9881, ZN => n1890);
   U8019 : OAI22_X1 port map( A1 => n10140, A2 => n9885, B1 => n7230, B2 => 
                           n9881, ZN => n1891);
   U8020 : OAI22_X1 port map( A1 => n10143, A2 => n9885, B1 => n7229, B2 => 
                           n9881, ZN => n1892);
   U8021 : OAI22_X1 port map( A1 => n10146, A2 => n9885, B1 => n7228, B2 => 
                           n9881, ZN => n1893);
   U8022 : OAI22_X1 port map( A1 => n10149, A2 => n9885, B1 => n7227, B2 => 
                           n9881, ZN => n1894);
   U8023 : OAI22_X1 port map( A1 => n10152, A2 => n9885, B1 => n7226, B2 => 
                           n9881, ZN => n1895);
   U8024 : OAI22_X1 port map( A1 => n10155, A2 => n9885, B1 => n7225, B2 => 
                           n9881, ZN => n1896);
   U8025 : OAI22_X1 port map( A1 => n10158, A2 => n9885, B1 => n7224, B2 => 
                           n9881, ZN => n1897);
   U8026 : OAI22_X1 port map( A1 => n10161, A2 => n9885, B1 => n7223, B2 => 
                           n9881, ZN => n1898);
   U8027 : OAI22_X1 port map( A1 => n10164, A2 => n9886, B1 => n7222, B2 => 
                           n9881, ZN => n1899);
   U8028 : OAI22_X1 port map( A1 => n10167, A2 => n9886, B1 => n7221, B2 => 
                           n9882, ZN => n1900);
   U8029 : OAI22_X1 port map( A1 => n10170, A2 => n9886, B1 => n7220, B2 => 
                           n9882, ZN => n1901);
   U8030 : OAI22_X1 port map( A1 => n10173, A2 => n9886, B1 => n7219, B2 => 
                           n9882, ZN => n1902);
   U8031 : OAI22_X1 port map( A1 => n10176, A2 => n9886, B1 => n7218, B2 => 
                           n9882, ZN => n1903);
   U8032 : OAI22_X1 port map( A1 => n10179, A2 => n9886, B1 => n7217, B2 => 
                           n9882, ZN => n1904);
   U8033 : OAI22_X1 port map( A1 => n10182, A2 => n9886, B1 => n7216, B2 => 
                           n9882, ZN => n1905);
   U8034 : OAI22_X1 port map( A1 => n10185, A2 => n9886, B1 => n7215, B2 => 
                           n9882, ZN => n1906);
   U8035 : OAI22_X1 port map( A1 => n10188, A2 => n9886, B1 => n7214, B2 => 
                           n9882, ZN => n1907);
   U8036 : OAI22_X1 port map( A1 => n10191, A2 => n9886, B1 => n7213, B2 => 
                           n9882, ZN => n1908);
   U8037 : OAI22_X1 port map( A1 => n10194, A2 => n9886, B1 => n7212, B2 => 
                           n9882, ZN => n1909);
   U8038 : OAI22_X1 port map( A1 => n10197, A2 => n9886, B1 => n7211, B2 => 
                           n9882, ZN => n1910);
   U8039 : OAI22_X1 port map( A1 => n10200, A2 => n9887, B1 => n7210, B2 => 
                           n9882, ZN => n1911);
   U8040 : OAI22_X1 port map( A1 => n10203, A2 => n9887, B1 => n7209, B2 => 
                           n9883, ZN => n1912);
   U8041 : OAI22_X1 port map( A1 => n10206, A2 => n9887, B1 => n7208, B2 => 
                           n9883, ZN => n1913);
   U8042 : OAI22_X1 port map( A1 => n10209, A2 => n9887, B1 => n7207, B2 => 
                           n9883, ZN => n1914);
   U8043 : OAI22_X1 port map( A1 => n10212, A2 => n9887, B1 => n7206, B2 => 
                           n9883, ZN => n1915);
   U8044 : OAI22_X1 port map( A1 => n10215, A2 => n9887, B1 => n7205, B2 => 
                           n9883, ZN => n1916);
   U8045 : OAI22_X1 port map( A1 => n10218, A2 => n9887, B1 => n7204, B2 => 
                           n9883, ZN => n1917);
   U8046 : OAI22_X1 port map( A1 => n10221, A2 => n9887, B1 => n7203, B2 => 
                           n9883, ZN => n1918);
   U8047 : OAI22_X1 port map( A1 => n10224, A2 => n9887, B1 => n7202, B2 => 
                           n9883, ZN => n1919);
   U8048 : OAI22_X1 port map( A1 => n10133, A2 => n9941, B1 => n7008, B2 => 
                           n9937, ZN => n2113);
   U8049 : OAI22_X1 port map( A1 => n10136, A2 => n9941, B1 => n7007, B2 => 
                           n9937, ZN => n2114);
   U8050 : OAI22_X1 port map( A1 => n10139, A2 => n9941, B1 => n7006, B2 => 
                           n9937, ZN => n2115);
   U8051 : OAI22_X1 port map( A1 => n10151, A2 => n9941, B1 => n7002, B2 => 
                           n9937, ZN => n2119);
   U8052 : OAI22_X1 port map( A1 => n10154, A2 => n9941, B1 => n7001, B2 => 
                           n9937, ZN => n2120);
   U8053 : OAI22_X1 port map( A1 => n10166, A2 => n9942, B1 => n6997, B2 => 
                           n9938, ZN => n2124);
   U8054 : OAI22_X1 port map( A1 => n10172, A2 => n9942, B1 => n6995, B2 => 
                           n9938, ZN => n2126);
   U8055 : OAI22_X1 port map( A1 => n10175, A2 => n9942, B1 => n6994, B2 => 
                           n9938, ZN => n2127);
   U8056 : OAI22_X1 port map( A1 => n10178, A2 => n9942, B1 => n6993, B2 => 
                           n9938, ZN => n2128);
   U8057 : OAI22_X1 port map( A1 => n10181, A2 => n9942, B1 => n6992, B2 => 
                           n9938, ZN => n2129);
   U8058 : OAI22_X1 port map( A1 => n10187, A2 => n9942, B1 => n6990, B2 => 
                           n9938, ZN => n2131);
   U8059 : OAI22_X1 port map( A1 => n10190, A2 => n9942, B1 => n6989, B2 => 
                           n9938, ZN => n2132);
   U8060 : OAI22_X1 port map( A1 => n10193, A2 => n9942, B1 => n6988, B2 => 
                           n9938, ZN => n2133);
   U8061 : OAI22_X1 port map( A1 => n10196, A2 => n9942, B1 => n6987, B2 => 
                           n9938, ZN => n2134);
   U8062 : OAI22_X1 port map( A1 => n10199, A2 => n9943, B1 => n6986, B2 => 
                           n9938, ZN => n2135);
   U8063 : OAI22_X1 port map( A1 => n10202, A2 => n9943, B1 => n6985, B2 => 
                           n9939, ZN => n2136);
   U8064 : OAI22_X1 port map( A1 => n10205, A2 => n9943, B1 => n6984, B2 => 
                           n9939, ZN => n2137);
   U8065 : OAI22_X1 port map( A1 => n10208, A2 => n9943, B1 => n6983, B2 => 
                           n9939, ZN => n2138);
   U8066 : OAI22_X1 port map( A1 => n10132, A2 => n9773, B1 => n7424, B2 => 
                           n9769, ZN => n1440);
   U8067 : OAI22_X1 port map( A1 => n10135, A2 => n9773, B1 => n7423, B2 => 
                           n9769, ZN => n1441);
   U8068 : OAI22_X1 port map( A1 => n10138, A2 => n9773, B1 => n7422, B2 => 
                           n9769, ZN => n1442);
   U8069 : OAI22_X1 port map( A1 => n10141, A2 => n9773, B1 => n7421, B2 => 
                           n9769, ZN => n1443);
   U8070 : OAI22_X1 port map( A1 => n10144, A2 => n9773, B1 => n7420, B2 => 
                           n9769, ZN => n1444);
   U8071 : OAI22_X1 port map( A1 => n10147, A2 => n9773, B1 => n7419, B2 => 
                           n9769, ZN => n1445);
   U8072 : OAI22_X1 port map( A1 => n10150, A2 => n9773, B1 => n7418, B2 => 
                           n9769, ZN => n1446);
   U8073 : OAI22_X1 port map( A1 => n10153, A2 => n9773, B1 => n7417, B2 => 
                           n9769, ZN => n1447);
   U8074 : OAI22_X1 port map( A1 => n10156, A2 => n9773, B1 => n7416, B2 => 
                           n9769, ZN => n1448);
   U8075 : OAI22_X1 port map( A1 => n10159, A2 => n9773, B1 => n7415, B2 => 
                           n9769, ZN => n1449);
   U8076 : OAI22_X1 port map( A1 => n10162, A2 => n9773, B1 => n7414, B2 => 
                           n9769, ZN => n1450);
   U8077 : OAI22_X1 port map( A1 => n10165, A2 => n9774, B1 => n7413, B2 => 
                           n9769, ZN => n1451);
   U8078 : OAI22_X1 port map( A1 => n10168, A2 => n9774, B1 => n7412, B2 => 
                           n9770, ZN => n1452);
   U8079 : OAI22_X1 port map( A1 => n10171, A2 => n9774, B1 => n7411, B2 => 
                           n9770, ZN => n1453);
   U8080 : OAI22_X1 port map( A1 => n10174, A2 => n9774, B1 => n7410, B2 => 
                           n9770, ZN => n1454);
   U8081 : OAI22_X1 port map( A1 => n10177, A2 => n9774, B1 => n7409, B2 => 
                           n9770, ZN => n1455);
   U8082 : OAI22_X1 port map( A1 => n10180, A2 => n9774, B1 => n7408, B2 => 
                           n9770, ZN => n1456);
   U8083 : OAI22_X1 port map( A1 => n10183, A2 => n9774, B1 => n7407, B2 => 
                           n9770, ZN => n1457);
   U8084 : OAI22_X1 port map( A1 => n10186, A2 => n9774, B1 => n7406, B2 => 
                           n9770, ZN => n1458);
   U8085 : OAI22_X1 port map( A1 => n10189, A2 => n9774, B1 => n7405, B2 => 
                           n9770, ZN => n1459);
   U8086 : OAI22_X1 port map( A1 => n10192, A2 => n9774, B1 => n7404, B2 => 
                           n9770, ZN => n1460);
   U8087 : OAI22_X1 port map( A1 => n10195, A2 => n9774, B1 => n7403, B2 => 
                           n9770, ZN => n1461);
   U8088 : OAI22_X1 port map( A1 => n10198, A2 => n9774, B1 => n7402, B2 => 
                           n9770, ZN => n1462);
   U8089 : OAI22_X1 port map( A1 => n10201, A2 => n9775, B1 => n7401, B2 => 
                           n9770, ZN => n1463);
   U8090 : OAI22_X1 port map( A1 => n10204, A2 => n9775, B1 => n7400, B2 => 
                           n9771, ZN => n1464);
   U8091 : OAI22_X1 port map( A1 => n10207, A2 => n9775, B1 => n7399, B2 => 
                           n9771, ZN => n1465);
   U8092 : OAI22_X1 port map( A1 => n10210, A2 => n9775, B1 => n7398, B2 => 
                           n9771, ZN => n1466);
   U8093 : OAI22_X1 port map( A1 => n10213, A2 => n9775, B1 => n7397, B2 => 
                           n9771, ZN => n1467);
   U8094 : OAI22_X1 port map( A1 => n10216, A2 => n9775, B1 => n7396, B2 => 
                           n9771, ZN => n1468);
   U8095 : OAI22_X1 port map( A1 => n10222, A2 => n9775, B1 => n7394, B2 => 
                           n9771, ZN => n1470);
   U8096 : OAI22_X1 port map( A1 => n10225, A2 => n9775, B1 => n7393, B2 => 
                           n9771, ZN => n1471);
   U8097 : OAI22_X1 port map( A1 => n10131, A2 => n9789, B1 => n7392, B2 => 
                           n9785, ZN => n1504);
   U8098 : OAI22_X1 port map( A1 => n10134, A2 => n9789, B1 => n7391, B2 => 
                           n9785, ZN => n1505);
   U8099 : OAI22_X1 port map( A1 => n10137, A2 => n9789, B1 => n7390, B2 => 
                           n9785, ZN => n1506);
   U8100 : OAI22_X1 port map( A1 => n10140, A2 => n9789, B1 => n7389, B2 => 
                           n9785, ZN => n1507);
   U8101 : OAI22_X1 port map( A1 => n10143, A2 => n9789, B1 => n7388, B2 => 
                           n9785, ZN => n1508);
   U8102 : OAI22_X1 port map( A1 => n10146, A2 => n9789, B1 => n7387, B2 => 
                           n9785, ZN => n1509);
   U8103 : OAI22_X1 port map( A1 => n10149, A2 => n9789, B1 => n7386, B2 => 
                           n9785, ZN => n1510);
   U8104 : OAI22_X1 port map( A1 => n10152, A2 => n9789, B1 => n7385, B2 => 
                           n9785, ZN => n1511);
   U8105 : OAI22_X1 port map( A1 => n10155, A2 => n9789, B1 => n7384, B2 => 
                           n9785, ZN => n1512);
   U8106 : OAI22_X1 port map( A1 => n10158, A2 => n9789, B1 => n7383, B2 => 
                           n9785, ZN => n1513);
   U8107 : OAI22_X1 port map( A1 => n10161, A2 => n9789, B1 => n7382, B2 => 
                           n9785, ZN => n1514);
   U8108 : OAI22_X1 port map( A1 => n10164, A2 => n9790, B1 => n7381, B2 => 
                           n9785, ZN => n1515);
   U8109 : OAI22_X1 port map( A1 => n10167, A2 => n9790, B1 => n7380, B2 => 
                           n9786, ZN => n1516);
   U8110 : OAI22_X1 port map( A1 => n10170, A2 => n9790, B1 => n7379, B2 => 
                           n9786, ZN => n1517);
   U8111 : OAI22_X1 port map( A1 => n10173, A2 => n9790, B1 => n7378, B2 => 
                           n9786, ZN => n1518);
   U8112 : OAI22_X1 port map( A1 => n10176, A2 => n9790, B1 => n7377, B2 => 
                           n9786, ZN => n1519);
   U8113 : OAI22_X1 port map( A1 => n10179, A2 => n9790, B1 => n7376, B2 => 
                           n9786, ZN => n1520);
   U8114 : OAI22_X1 port map( A1 => n10182, A2 => n9790, B1 => n7375, B2 => 
                           n9786, ZN => n1521);
   U8115 : OAI22_X1 port map( A1 => n10185, A2 => n9790, B1 => n7374, B2 => 
                           n9786, ZN => n1522);
   U8116 : OAI22_X1 port map( A1 => n10188, A2 => n9790, B1 => n7373, B2 => 
                           n9786, ZN => n1523);
   U8117 : OAI22_X1 port map( A1 => n10191, A2 => n9790, B1 => n7372, B2 => 
                           n9786, ZN => n1524);
   U8118 : OAI22_X1 port map( A1 => n10194, A2 => n9790, B1 => n7371, B2 => 
                           n9786, ZN => n1525);
   U8119 : OAI22_X1 port map( A1 => n10197, A2 => n9790, B1 => n7370, B2 => 
                           n9786, ZN => n1526);
   U8120 : OAI22_X1 port map( A1 => n10200, A2 => n9791, B1 => n7369, B2 => 
                           n9786, ZN => n1527);
   U8121 : OAI22_X1 port map( A1 => n10203, A2 => n9791, B1 => n7368, B2 => 
                           n9787, ZN => n1528);
   U8122 : OAI22_X1 port map( A1 => n10206, A2 => n9791, B1 => n7367, B2 => 
                           n9787, ZN => n1529);
   U8123 : OAI22_X1 port map( A1 => n10209, A2 => n9791, B1 => n7366, B2 => 
                           n9787, ZN => n1530);
   U8124 : OAI22_X1 port map( A1 => n10218, A2 => n9791, B1 => n7363, B2 => 
                           n9787, ZN => n1533);
   U8125 : OAI22_X1 port map( A1 => n10224, A2 => n9791, B1 => n7361, B2 => 
                           n9787, ZN => n1535);
   U8126 : OAI22_X1 port map( A1 => n10131, A2 => n9837, B1 => n7360, B2 => 
                           n9833, ZN => n1696);
   U8127 : OAI22_X1 port map( A1 => n10134, A2 => n9837, B1 => n7359, B2 => 
                           n9833, ZN => n1697);
   U8128 : OAI22_X1 port map( A1 => n10137, A2 => n9837, B1 => n7358, B2 => 
                           n9833, ZN => n1698);
   U8129 : OAI22_X1 port map( A1 => n10140, A2 => n9837, B1 => n7357, B2 => 
                           n9833, ZN => n1699);
   U8130 : OAI22_X1 port map( A1 => n10143, A2 => n9837, B1 => n7356, B2 => 
                           n9833, ZN => n1700);
   U8131 : OAI22_X1 port map( A1 => n10146, A2 => n9837, B1 => n7355, B2 => 
                           n9833, ZN => n1701);
   U8132 : OAI22_X1 port map( A1 => n10149, A2 => n9837, B1 => n7354, B2 => 
                           n9833, ZN => n1702);
   U8133 : OAI22_X1 port map( A1 => n10152, A2 => n9837, B1 => n7353, B2 => 
                           n9833, ZN => n1703);
   U8134 : OAI22_X1 port map( A1 => n10155, A2 => n9837, B1 => n7352, B2 => 
                           n9833, ZN => n1704);
   U8135 : OAI22_X1 port map( A1 => n10158, A2 => n9837, B1 => n7351, B2 => 
                           n9833, ZN => n1705);
   U8136 : OAI22_X1 port map( A1 => n10161, A2 => n9837, B1 => n7350, B2 => 
                           n9833, ZN => n1706);
   U8137 : OAI22_X1 port map( A1 => n10164, A2 => n9838, B1 => n7349, B2 => 
                           n9833, ZN => n1707);
   U8138 : OAI22_X1 port map( A1 => n10167, A2 => n9838, B1 => n7348, B2 => 
                           n9834, ZN => n1708);
   U8139 : OAI22_X1 port map( A1 => n10173, A2 => n9838, B1 => n7346, B2 => 
                           n9834, ZN => n1710);
   U8140 : OAI22_X1 port map( A1 => n10176, A2 => n9838, B1 => n7345, B2 => 
                           n9834, ZN => n1711);
   U8141 : OAI22_X1 port map( A1 => n10179, A2 => n9838, B1 => n7344, B2 => 
                           n9834, ZN => n1712);
   U8142 : OAI22_X1 port map( A1 => n10182, A2 => n9838, B1 => n7343, B2 => 
                           n9834, ZN => n1713);
   U8143 : OAI22_X1 port map( A1 => n10185, A2 => n9838, B1 => n7342, B2 => 
                           n9834, ZN => n1714);
   U8144 : OAI22_X1 port map( A1 => n10191, A2 => n9838, B1 => n7340, B2 => 
                           n9834, ZN => n1716);
   U8145 : OAI22_X1 port map( A1 => n10194, A2 => n9838, B1 => n7339, B2 => 
                           n9834, ZN => n1717);
   U8146 : OAI22_X1 port map( A1 => n10197, A2 => n9838, B1 => n7338, B2 => 
                           n9834, ZN => n1718);
   U8147 : OAI22_X1 port map( A1 => n10200, A2 => n9839, B1 => n7337, B2 => 
                           n9834, ZN => n1719);
   U8148 : OAI22_X1 port map( A1 => n10203, A2 => n9839, B1 => n7336, B2 => 
                           n9835, ZN => n1720);
   U8149 : OAI22_X1 port map( A1 => n10206, A2 => n9839, B1 => n7335, B2 => 
                           n9835, ZN => n1721);
   U8150 : OAI22_X1 port map( A1 => n10209, A2 => n9839, B1 => n7334, B2 => 
                           n9835, ZN => n1722);
   U8151 : OAI22_X1 port map( A1 => n10212, A2 => n9839, B1 => n7333, B2 => 
                           n9835, ZN => n1723);
   U8152 : OAI22_X1 port map( A1 => n10215, A2 => n9839, B1 => n7332, B2 => 
                           n9835, ZN => n1724);
   U8153 : OAI22_X1 port map( A1 => n10218, A2 => n9839, B1 => n7331, B2 => 
                           n9835, ZN => n1725);
   U8154 : OAI22_X1 port map( A1 => n10221, A2 => n9839, B1 => n7330, B2 => 
                           n9835, ZN => n1726);
   U8155 : OAI22_X1 port map( A1 => n10224, A2 => n9839, B1 => n7329, B2 => 
                           n9835, ZN => n1727);
   U8156 : OAI22_X1 port map( A1 => n10134, A2 => n9877, B1 => n7264, B2 => 
                           n9873, ZN => n1857);
   U8157 : OAI22_X1 port map( A1 => n10137, A2 => n9877, B1 => n7263, B2 => 
                           n9873, ZN => n1858);
   U8158 : OAI22_X1 port map( A1 => n10140, A2 => n9877, B1 => n7262, B2 => 
                           n9873, ZN => n1859);
   U8159 : OAI22_X1 port map( A1 => n10143, A2 => n9877, B1 => n7261, B2 => 
                           n9873, ZN => n1860);
   U8160 : OAI22_X1 port map( A1 => n10146, A2 => n9877, B1 => n7260, B2 => 
                           n9873, ZN => n1861);
   U8161 : OAI22_X1 port map( A1 => n10149, A2 => n9877, B1 => n7259, B2 => 
                           n9873, ZN => n1862);
   U8162 : OAI22_X1 port map( A1 => n10152, A2 => n9877, B1 => n7258, B2 => 
                           n9873, ZN => n1863);
   U8163 : OAI22_X1 port map( A1 => n10155, A2 => n9877, B1 => n7257, B2 => 
                           n9873, ZN => n1864);
   U8164 : OAI22_X1 port map( A1 => n10158, A2 => n9877, B1 => n7256, B2 => 
                           n9873, ZN => n1865);
   U8165 : OAI22_X1 port map( A1 => n10161, A2 => n9877, B1 => n7255, B2 => 
                           n9873, ZN => n1866);
   U8166 : OAI22_X1 port map( A1 => n10170, A2 => n9878, B1 => n7252, B2 => 
                           n9874, ZN => n1869);
   U8167 : OAI22_X1 port map( A1 => n10173, A2 => n9878, B1 => n7251, B2 => 
                           n9874, ZN => n1870);
   U8168 : OAI22_X1 port map( A1 => n10176, A2 => n9878, B1 => n7250, B2 => 
                           n9874, ZN => n1871);
   U8169 : OAI22_X1 port map( A1 => n10179, A2 => n9878, B1 => n7249, B2 => 
                           n9874, ZN => n1872);
   U8170 : OAI22_X1 port map( A1 => n10182, A2 => n9878, B1 => n7248, B2 => 
                           n9874, ZN => n1873);
   U8171 : OAI22_X1 port map( A1 => n10188, A2 => n9878, B1 => n7246, B2 => 
                           n9874, ZN => n1875);
   U8172 : OAI22_X1 port map( A1 => n10191, A2 => n9878, B1 => n7245, B2 => 
                           n9874, ZN => n1876);
   U8173 : OAI22_X1 port map( A1 => n10194, A2 => n9878, B1 => n7244, B2 => 
                           n9874, ZN => n1877);
   U8174 : OAI22_X1 port map( A1 => n10197, A2 => n9878, B1 => n7243, B2 => 
                           n9874, ZN => n1878);
   U8175 : OAI22_X1 port map( A1 => n10200, A2 => n9879, B1 => n7242, B2 => 
                           n9874, ZN => n1879);
   U8176 : OAI22_X1 port map( A1 => n10203, A2 => n9879, B1 => n7241, B2 => 
                           n9875, ZN => n1880);
   U8177 : OAI22_X1 port map( A1 => n10206, A2 => n9879, B1 => n7240, B2 => 
                           n9875, ZN => n1881);
   U8178 : OAI22_X1 port map( A1 => n10209, A2 => n9879, B1 => n7239, B2 => 
                           n9875, ZN => n1882);
   U8179 : OAI22_X1 port map( A1 => n10212, A2 => n9879, B1 => n7238, B2 => 
                           n9875, ZN => n1883);
   U8180 : OAI22_X1 port map( A1 => n10215, A2 => n9879, B1 => n7237, B2 => 
                           n9875, ZN => n1884);
   U8181 : OAI22_X1 port map( A1 => n10218, A2 => n9879, B1 => n7236, B2 => 
                           n9875, ZN => n1885);
   U8182 : OAI22_X1 port map( A1 => n10221, A2 => n9879, B1 => n7235, B2 => 
                           n9875, ZN => n1886);
   U8183 : OAI22_X1 port map( A1 => n10224, A2 => n9879, B1 => n7234, B2 => 
                           n9875, ZN => n1887);
   U8184 : OAI22_X1 port map( A1 => n10130, A2 => n9909, B1 => n7137, B2 => 
                           n9905, ZN => n1984);
   U8185 : OAI22_X1 port map( A1 => n10139, A2 => n9909, B1 => n7134, B2 => 
                           n9905, ZN => n1987);
   U8186 : OAI22_X1 port map( A1 => n10142, A2 => n9909, B1 => n7133, B2 => 
                           n9905, ZN => n1988);
   U8187 : OAI22_X1 port map( A1 => n10145, A2 => n9909, B1 => n7132, B2 => 
                           n9905, ZN => n1989);
   U8188 : OAI22_X1 port map( A1 => n10148, A2 => n9909, B1 => n7131, B2 => 
                           n9905, ZN => n1990);
   U8189 : OAI22_X1 port map( A1 => n10151, A2 => n9909, B1 => n7130, B2 => 
                           n9905, ZN => n1991);
   U8190 : OAI22_X1 port map( A1 => n10154, A2 => n9909, B1 => n7129, B2 => 
                           n9905, ZN => n1992);
   U8191 : OAI22_X1 port map( A1 => n10157, A2 => n9909, B1 => n7128, B2 => 
                           n9905, ZN => n1993);
   U8192 : OAI22_X1 port map( A1 => n10160, A2 => n9909, B1 => n7127, B2 => 
                           n9905, ZN => n1994);
   U8193 : OAI22_X1 port map( A1 => n10166, A2 => n9910, B1 => n7125, B2 => 
                           n9906, ZN => n1996);
   U8194 : OAI22_X1 port map( A1 => n10169, A2 => n9910, B1 => n7124, B2 => 
                           n9906, ZN => n1997);
   U8195 : OAI22_X1 port map( A1 => n10172, A2 => n9910, B1 => n7123, B2 => 
                           n9906, ZN => n1998);
   U8196 : OAI22_X1 port map( A1 => n10175, A2 => n9910, B1 => n7122, B2 => 
                           n9906, ZN => n1999);
   U8197 : OAI22_X1 port map( A1 => n10178, A2 => n9910, B1 => n7121, B2 => 
                           n9906, ZN => n2000);
   U8198 : OAI22_X1 port map( A1 => n10181, A2 => n9910, B1 => n7120, B2 => 
                           n9906, ZN => n2001);
   U8199 : OAI22_X1 port map( A1 => n10184, A2 => n9910, B1 => n7119, B2 => 
                           n9906, ZN => n2002);
   U8200 : OAI22_X1 port map( A1 => n10187, A2 => n9910, B1 => n7118, B2 => 
                           n9906, ZN => n2003);
   U8201 : OAI22_X1 port map( A1 => n10190, A2 => n9910, B1 => n7117, B2 => 
                           n9906, ZN => n2004);
   U8202 : OAI22_X1 port map( A1 => n10193, A2 => n9910, B1 => n7116, B2 => 
                           n9906, ZN => n2005);
   U8203 : OAI22_X1 port map( A1 => n10196, A2 => n9910, B1 => n7115, B2 => 
                           n9906, ZN => n2006);
   U8204 : OAI22_X1 port map( A1 => n10199, A2 => n9911, B1 => n7114, B2 => 
                           n9906, ZN => n2007);
   U8205 : OAI22_X1 port map( A1 => n10202, A2 => n9911, B1 => n7113, B2 => 
                           n9907, ZN => n2008);
   U8206 : OAI22_X1 port map( A1 => n10205, A2 => n9911, B1 => n7112, B2 => 
                           n9907, ZN => n2009);
   U8207 : OAI22_X1 port map( A1 => n10208, A2 => n9911, B1 => n7111, B2 => 
                           n9907, ZN => n2010);
   U8208 : OAI22_X1 port map( A1 => n10211, A2 => n9911, B1 => n7110, B2 => 
                           n9907, ZN => n2011);
   U8209 : OAI22_X1 port map( A1 => n10214, A2 => n9911, B1 => n7109, B2 => 
                           n9907, ZN => n2012);
   U8210 : OAI22_X1 port map( A1 => n10217, A2 => n9911, B1 => n7108, B2 => 
                           n9907, ZN => n2013);
   U8211 : OAI22_X1 port map( A1 => n10220, A2 => n9911, B1 => n7107, B2 => 
                           n9907, ZN => n2014);
   U8212 : OAI22_X1 port map( A1 => n10223, A2 => n9911, B1 => n7106, B2 => 
                           n9907, ZN => n2015);
   U8213 : OAI22_X1 port map( A1 => n10130, A2 => n9941, B1 => n7009, B2 => 
                           n9937, ZN => n2112);
   U8214 : OAI22_X1 port map( A1 => n10142, A2 => n9941, B1 => n7005, B2 => 
                           n9937, ZN => n2116);
   U8215 : OAI22_X1 port map( A1 => n10145, A2 => n9941, B1 => n7004, B2 => 
                           n9937, ZN => n2117);
   U8216 : OAI22_X1 port map( A1 => n10148, A2 => n9941, B1 => n7003, B2 => 
                           n9937, ZN => n2118);
   U8217 : OAI22_X1 port map( A1 => n10157, A2 => n9941, B1 => n7000, B2 => 
                           n9937, ZN => n2121);
   U8218 : OAI22_X1 port map( A1 => n10160, A2 => n9941, B1 => n6999, B2 => 
                           n9937, ZN => n2122);
   U8219 : OAI22_X1 port map( A1 => n10163, A2 => n9942, B1 => n6998, B2 => 
                           n9937, ZN => n2123);
   U8220 : OAI22_X1 port map( A1 => n10169, A2 => n9942, B1 => n6996, B2 => 
                           n9938, ZN => n2125);
   U8221 : OAI22_X1 port map( A1 => n10184, A2 => n9942, B1 => n6991, B2 => 
                           n9938, ZN => n2130);
   U8222 : OAI22_X1 port map( A1 => n10211, A2 => n9943, B1 => n6982, B2 => 
                           n9939, ZN => n2139);
   U8223 : OAI22_X1 port map( A1 => n10214, A2 => n9943, B1 => n6981, B2 => 
                           n9939, ZN => n2140);
   U8224 : OAI22_X1 port map( A1 => n10217, A2 => n9943, B1 => n6980, B2 => 
                           n9939, ZN => n2141);
   U8225 : OAI22_X1 port map( A1 => n10220, A2 => n9943, B1 => n6979, B2 => 
                           n9939, ZN => n2142);
   U8226 : OAI22_X1 port map( A1 => n10223, A2 => n9943, B1 => n6978, B2 => 
                           n9939, ZN => n2143);
   U8227 : OAI22_X1 port map( A1 => n10219, A2 => n9775, B1 => n7395, B2 => 
                           n9771, ZN => n1469);
   U8228 : OAI22_X1 port map( A1 => n10212, A2 => n9791, B1 => n7365, B2 => 
                           n9787, ZN => n1531);
   U8229 : OAI22_X1 port map( A1 => n10215, A2 => n9791, B1 => n7364, B2 => 
                           n9787, ZN => n1532);
   U8230 : OAI22_X1 port map( A1 => n10221, A2 => n9791, B1 => n7362, B2 => 
                           n9787, ZN => n1534);
   U8231 : OAI22_X1 port map( A1 => n10170, A2 => n9838, B1 => n7347, B2 => 
                           n9834, ZN => n1709);
   U8232 : OAI22_X1 port map( A1 => n10188, A2 => n9838, B1 => n7341, B2 => 
                           n9834, ZN => n1715);
   U8233 : OAI22_X1 port map( A1 => n10131, A2 => n9877, B1 => n7265, B2 => 
                           n9873, ZN => n1856);
   U8234 : OAI22_X1 port map( A1 => n10164, A2 => n9878, B1 => n7254, B2 => 
                           n9873, ZN => n1867);
   U8235 : OAI22_X1 port map( A1 => n10167, A2 => n9878, B1 => n7253, B2 => 
                           n9874, ZN => n1868);
   U8236 : OAI22_X1 port map( A1 => n10185, A2 => n9878, B1 => n7247, B2 => 
                           n9874, ZN => n1874);
   U8237 : OAI22_X1 port map( A1 => n10133, A2 => n9909, B1 => n7136, B2 => 
                           n9905, ZN => n1985);
   U8238 : OAI22_X1 port map( A1 => n10136, A2 => n9909, B1 => n7135, B2 => 
                           n9905, ZN => n1986);
   U8239 : OAI22_X1 port map( A1 => n10163, A2 => n9910, B1 => n7126, B2 => 
                           n9905, ZN => n1995);
   U8240 : OAI22_X1 port map( A1 => n10130, A2 => n9917, B1 => n7105, B2 => 
                           n9913, ZN => n2016);
   U8241 : OAI22_X1 port map( A1 => n10133, A2 => n9917, B1 => n7104, B2 => 
                           n9913, ZN => n2017);
   U8242 : OAI22_X1 port map( A1 => n10136, A2 => n9917, B1 => n7103, B2 => 
                           n9913, ZN => n2018);
   U8243 : OAI22_X1 port map( A1 => n10139, A2 => n9917, B1 => n7102, B2 => 
                           n9913, ZN => n2019);
   U8244 : OAI22_X1 port map( A1 => n10142, A2 => n9917, B1 => n7101, B2 => 
                           n9913, ZN => n2020);
   U8245 : OAI22_X1 port map( A1 => n10145, A2 => n9917, B1 => n7100, B2 => 
                           n9913, ZN => n2021);
   U8246 : OAI22_X1 port map( A1 => n10148, A2 => n9917, B1 => n7099, B2 => 
                           n9913, ZN => n2022);
   U8247 : OAI22_X1 port map( A1 => n10151, A2 => n9917, B1 => n7098, B2 => 
                           n9913, ZN => n2023);
   U8248 : OAI22_X1 port map( A1 => n10154, A2 => n9917, B1 => n7097, B2 => 
                           n9913, ZN => n2024);
   U8249 : OAI22_X1 port map( A1 => n10157, A2 => n9917, B1 => n7096, B2 => 
                           n9913, ZN => n2025);
   U8250 : OAI22_X1 port map( A1 => n10160, A2 => n9917, B1 => n7095, B2 => 
                           n9913, ZN => n2026);
   U8251 : OAI22_X1 port map( A1 => n10163, A2 => n9918, B1 => n7094, B2 => 
                           n9913, ZN => n2027);
   U8252 : OAI22_X1 port map( A1 => n10166, A2 => n9918, B1 => n7093, B2 => 
                           n9914, ZN => n2028);
   U8253 : OAI22_X1 port map( A1 => n10169, A2 => n9918, B1 => n7092, B2 => 
                           n9914, ZN => n2029);
   U8254 : OAI22_X1 port map( A1 => n10172, A2 => n9918, B1 => n7091, B2 => 
                           n9914, ZN => n2030);
   U8255 : OAI22_X1 port map( A1 => n10175, A2 => n9918, B1 => n7090, B2 => 
                           n9914, ZN => n2031);
   U8256 : OAI22_X1 port map( A1 => n10178, A2 => n9918, B1 => n7089, B2 => 
                           n9914, ZN => n2032);
   U8257 : OAI22_X1 port map( A1 => n10181, A2 => n9918, B1 => n7088, B2 => 
                           n9914, ZN => n2033);
   U8258 : OAI22_X1 port map( A1 => n10184, A2 => n9918, B1 => n7087, B2 => 
                           n9914, ZN => n2034);
   U8259 : OAI22_X1 port map( A1 => n10187, A2 => n9918, B1 => n7086, B2 => 
                           n9914, ZN => n2035);
   U8260 : OAI22_X1 port map( A1 => n10190, A2 => n9918, B1 => n7085, B2 => 
                           n9914, ZN => n2036);
   U8261 : OAI22_X1 port map( A1 => n10193, A2 => n9918, B1 => n7084, B2 => 
                           n9914, ZN => n2037);
   U8262 : OAI22_X1 port map( A1 => n10196, A2 => n9918, B1 => n7083, B2 => 
                           n9914, ZN => n2038);
   U8263 : OAI22_X1 port map( A1 => n10199, A2 => n9919, B1 => n7082, B2 => 
                           n9914, ZN => n2039);
   U8264 : OAI22_X1 port map( A1 => n10202, A2 => n9919, B1 => n7081, B2 => 
                           n9915, ZN => n2040);
   U8265 : OAI22_X1 port map( A1 => n10205, A2 => n9919, B1 => n7080, B2 => 
                           n9915, ZN => n2041);
   U8266 : OAI22_X1 port map( A1 => n10208, A2 => n9919, B1 => n7079, B2 => 
                           n9915, ZN => n2042);
   U8267 : OAI22_X1 port map( A1 => n10211, A2 => n9919, B1 => n7078, B2 => 
                           n9915, ZN => n2043);
   U8268 : OAI22_X1 port map( A1 => n10214, A2 => n9919, B1 => n7077, B2 => 
                           n9915, ZN => n2044);
   U8269 : OAI22_X1 port map( A1 => n10217, A2 => n9919, B1 => n7076, B2 => 
                           n9915, ZN => n2045);
   U8270 : OAI22_X1 port map( A1 => n10220, A2 => n9919, B1 => n7075, B2 => 
                           n9915, ZN => n2046);
   U8271 : OAI22_X1 port map( A1 => n10223, A2 => n9919, B1 => n7074, B2 => 
                           n9915, ZN => n2047);
   U8272 : OAI22_X1 port map( A1 => n10130, A2 => n9933, B1 => n7041, B2 => 
                           n9929, ZN => n2080);
   U8273 : OAI22_X1 port map( A1 => n10133, A2 => n9933, B1 => n7040, B2 => 
                           n9929, ZN => n2081);
   U8274 : OAI22_X1 port map( A1 => n10136, A2 => n9933, B1 => n7039, B2 => 
                           n9929, ZN => n2082);
   U8275 : OAI22_X1 port map( A1 => n10139, A2 => n9933, B1 => n7038, B2 => 
                           n9929, ZN => n2083);
   U8276 : OAI22_X1 port map( A1 => n10142, A2 => n9933, B1 => n7037, B2 => 
                           n9929, ZN => n2084);
   U8277 : OAI22_X1 port map( A1 => n10145, A2 => n9933, B1 => n7036, B2 => 
                           n9929, ZN => n2085);
   U8278 : OAI22_X1 port map( A1 => n10148, A2 => n9933, B1 => n7035, B2 => 
                           n9929, ZN => n2086);
   U8279 : OAI22_X1 port map( A1 => n10151, A2 => n9933, B1 => n7034, B2 => 
                           n9929, ZN => n2087);
   U8280 : OAI22_X1 port map( A1 => n10154, A2 => n9933, B1 => n7033, B2 => 
                           n9929, ZN => n2088);
   U8281 : OAI22_X1 port map( A1 => n10157, A2 => n9933, B1 => n7032, B2 => 
                           n9929, ZN => n2089);
   U8282 : OAI22_X1 port map( A1 => n10160, A2 => n9933, B1 => n7031, B2 => 
                           n9929, ZN => n2090);
   U8283 : OAI22_X1 port map( A1 => n10163, A2 => n9934, B1 => n7030, B2 => 
                           n9929, ZN => n2091);
   U8284 : OAI22_X1 port map( A1 => n10166, A2 => n9934, B1 => n7029, B2 => 
                           n9930, ZN => n2092);
   U8285 : OAI22_X1 port map( A1 => n10169, A2 => n9934, B1 => n7028, B2 => 
                           n9930, ZN => n2093);
   U8286 : OAI22_X1 port map( A1 => n10172, A2 => n9934, B1 => n7027, B2 => 
                           n9930, ZN => n2094);
   U8287 : OAI22_X1 port map( A1 => n10175, A2 => n9934, B1 => n7026, B2 => 
                           n9930, ZN => n2095);
   U8288 : OAI22_X1 port map( A1 => n10178, A2 => n9934, B1 => n7025, B2 => 
                           n9930, ZN => n2096);
   U8289 : OAI22_X1 port map( A1 => n10181, A2 => n9934, B1 => n7024, B2 => 
                           n9930, ZN => n2097);
   U8290 : OAI22_X1 port map( A1 => n10184, A2 => n9934, B1 => n7023, B2 => 
                           n9930, ZN => n2098);
   U8291 : OAI22_X1 port map( A1 => n10187, A2 => n9934, B1 => n7022, B2 => 
                           n9930, ZN => n2099);
   U8292 : OAI22_X1 port map( A1 => n10190, A2 => n9934, B1 => n7021, B2 => 
                           n9930, ZN => n2100);
   U8293 : OAI22_X1 port map( A1 => n10193, A2 => n9934, B1 => n7020, B2 => 
                           n9930, ZN => n2101);
   U8294 : OAI22_X1 port map( A1 => n10196, A2 => n9934, B1 => n7019, B2 => 
                           n9930, ZN => n2102);
   U8295 : OAI22_X1 port map( A1 => n10199, A2 => n9935, B1 => n7018, B2 => 
                           n9930, ZN => n2103);
   U8296 : OAI22_X1 port map( A1 => n10202, A2 => n9935, B1 => n7017, B2 => 
                           n9931, ZN => n2104);
   U8297 : OAI22_X1 port map( A1 => n10205, A2 => n9935, B1 => n7016, B2 => 
                           n9931, ZN => n2105);
   U8298 : OAI22_X1 port map( A1 => n10208, A2 => n9935, B1 => n7015, B2 => 
                           n9931, ZN => n2106);
   U8299 : OAI22_X1 port map( A1 => n10211, A2 => n9935, B1 => n7014, B2 => 
                           n9931, ZN => n2107);
   U8300 : OAI22_X1 port map( A1 => n10214, A2 => n9935, B1 => n7013, B2 => 
                           n9931, ZN => n2108);
   U8301 : OAI22_X1 port map( A1 => n10217, A2 => n9935, B1 => n7012, B2 => 
                           n9931, ZN => n2109);
   U8302 : OAI22_X1 port map( A1 => n10220, A2 => n9935, B1 => n7011, B2 => 
                           n9931, ZN => n2110);
   U8303 : OAI22_X1 port map( A1 => n10223, A2 => n9935, B1 => n7010, B2 => 
                           n9931, ZN => n2111);
   U8304 : OAI22_X1 port map( A1 => n10130, A2 => n9949, B1 => n6977, B2 => 
                           n9945, ZN => n2144);
   U8305 : OAI22_X1 port map( A1 => n10133, A2 => n9949, B1 => n6976, B2 => 
                           n9945, ZN => n2145);
   U8306 : OAI22_X1 port map( A1 => n10136, A2 => n9949, B1 => n6975, B2 => 
                           n9945, ZN => n2146);
   U8307 : OAI22_X1 port map( A1 => n10139, A2 => n9949, B1 => n6974, B2 => 
                           n9945, ZN => n2147);
   U8308 : OAI22_X1 port map( A1 => n10142, A2 => n9949, B1 => n6973, B2 => 
                           n9945, ZN => n2148);
   U8309 : OAI22_X1 port map( A1 => n10145, A2 => n9949, B1 => n6972, B2 => 
                           n9945, ZN => n2149);
   U8310 : OAI22_X1 port map( A1 => n10148, A2 => n9949, B1 => n6971, B2 => 
                           n9945, ZN => n2150);
   U8311 : OAI22_X1 port map( A1 => n10151, A2 => n9949, B1 => n6970, B2 => 
                           n9945, ZN => n2151);
   U8312 : OAI22_X1 port map( A1 => n10154, A2 => n9949, B1 => n6969, B2 => 
                           n9945, ZN => n2152);
   U8313 : OAI22_X1 port map( A1 => n10157, A2 => n9949, B1 => n6968, B2 => 
                           n9945, ZN => n2153);
   U8314 : OAI22_X1 port map( A1 => n10160, A2 => n9949, B1 => n6967, B2 => 
                           n9945, ZN => n2154);
   U8315 : OAI22_X1 port map( A1 => n10163, A2 => n9950, B1 => n6966, B2 => 
                           n9945, ZN => n2155);
   U8316 : OAI22_X1 port map( A1 => n10166, A2 => n9950, B1 => n6965, B2 => 
                           n9946, ZN => n2156);
   U8317 : OAI22_X1 port map( A1 => n10169, A2 => n9950, B1 => n6964, B2 => 
                           n9946, ZN => n2157);
   U8318 : OAI22_X1 port map( A1 => n10172, A2 => n9950, B1 => n6963, B2 => 
                           n9946, ZN => n2158);
   U8319 : OAI22_X1 port map( A1 => n10175, A2 => n9950, B1 => n6962, B2 => 
                           n9946, ZN => n2159);
   U8320 : OAI22_X1 port map( A1 => n10178, A2 => n9950, B1 => n6961, B2 => 
                           n9946, ZN => n2160);
   U8321 : OAI22_X1 port map( A1 => n10181, A2 => n9950, B1 => n6960, B2 => 
                           n9946, ZN => n2161);
   U8322 : OAI22_X1 port map( A1 => n10184, A2 => n9950, B1 => n6959, B2 => 
                           n9946, ZN => n2162);
   U8323 : OAI22_X1 port map( A1 => n10187, A2 => n9950, B1 => n6958, B2 => 
                           n9946, ZN => n2163);
   U8324 : OAI22_X1 port map( A1 => n10190, A2 => n9950, B1 => n6957, B2 => 
                           n9946, ZN => n2164);
   U8325 : OAI22_X1 port map( A1 => n10193, A2 => n9950, B1 => n6956, B2 => 
                           n9946, ZN => n2165);
   U8326 : OAI22_X1 port map( A1 => n10196, A2 => n9950, B1 => n6955, B2 => 
                           n9946, ZN => n2166);
   U8327 : OAI22_X1 port map( A1 => n10199, A2 => n9951, B1 => n6954, B2 => 
                           n9946, ZN => n2167);
   U8328 : OAI22_X1 port map( A1 => n10202, A2 => n9951, B1 => n6953, B2 => 
                           n9947, ZN => n2168);
   U8329 : OAI22_X1 port map( A1 => n10205, A2 => n9951, B1 => n6952, B2 => 
                           n9947, ZN => n2169);
   U8330 : OAI22_X1 port map( A1 => n10208, A2 => n9951, B1 => n6951, B2 => 
                           n9947, ZN => n2170);
   U8331 : OAI22_X1 port map( A1 => n10211, A2 => n9951, B1 => n6950, B2 => 
                           n9947, ZN => n2171);
   U8332 : OAI22_X1 port map( A1 => n10214, A2 => n9951, B1 => n6949, B2 => 
                           n9947, ZN => n2172);
   U8333 : OAI22_X1 port map( A1 => n10217, A2 => n9951, B1 => n6948, B2 => 
                           n9947, ZN => n2173);
   U8334 : OAI22_X1 port map( A1 => n10220, A2 => n9951, B1 => n6947, B2 => 
                           n9947, ZN => n2174);
   U8335 : OAI22_X1 port map( A1 => n10223, A2 => n9951, B1 => n6946, B2 => 
                           n9947, ZN => n2175);
   U8336 : NOR3_X1 port map( A1 => n6747, A2 => n6748, A3 => n6749, ZN => n8877
                           );
   U8337 : NOR3_X1 port map( A1 => n6751, A2 => n6752, A3 => n6753, ZN => n8209
                           );
   U8338 : AND3_X1 port map( A1 => n6744, A2 => n6743, A3 => n8237, ZN => n8227
                           );
   U8339 : AND3_X1 port map( A1 => n6744, A2 => n6743, A3 => n8274, ZN => n8267
                           );
   U8340 : NAND2_X1 port map( A1 => n8887, A2 => n8877, ZN => n8336);
   U8341 : NAND2_X1 port map( A1 => n8887, A2 => n8878, ZN => n8335);
   U8342 : NAND2_X1 port map( A1 => n8888, A2 => n8878, ZN => n8334);
   U8343 : NAND2_X1 port map( A1 => n8888, A2 => n8869, ZN => n8347);
   U8344 : NAND2_X1 port map( A1 => n8888, A2 => n8875, ZN => n8346);
   U8345 : NAND2_X1 port map( A1 => n8887, A2 => n8869, ZN => n8345);
   U8346 : NAND2_X1 port map( A1 => n8887, A2 => n8870, ZN => n8340);
   U8347 : NAND2_X1 port map( A1 => n8888, A2 => n8871, ZN => n8341);
   U8348 : NAND2_X1 port map( A1 => n8877, A2 => n8868, ZN => n8351);
   U8349 : NAND2_X1 port map( A1 => n8878, A2 => n8868, ZN => n8352);
   U8350 : NAND2_X1 port map( A1 => n8219, A2 => n8209, ZN => n7668);
   U8351 : NAND2_X1 port map( A1 => n8219, A2 => n8210, ZN => n7667);
   U8352 : NAND2_X1 port map( A1 => n8220, A2 => n8210, ZN => n7666);
   U8353 : NAND2_X1 port map( A1 => n8220, A2 => n8201, ZN => n7679);
   U8354 : NAND2_X1 port map( A1 => n8220, A2 => n8207, ZN => n7678);
   U8355 : NAND2_X1 port map( A1 => n8219, A2 => n8201, ZN => n7677);
   U8356 : NAND2_X1 port map( A1 => n8220, A2 => n8203, ZN => n7673);
   U8357 : NAND2_X1 port map( A1 => n8219, A2 => n8202, ZN => n7672);
   U8358 : NAND2_X1 port map( A1 => n8209, A2 => n8200, ZN => n7683);
   U8359 : NAND2_X1 port map( A1 => n8210, A2 => n8200, ZN => n7684);
   U8360 : NAND2_X1 port map( A1 => n8267, A2 => n8226, ZN => n8265);
   U8361 : NAND2_X1 port map( A1 => n8267, A2 => n8233, ZN => n8270);
   U8362 : NAND2_X1 port map( A1 => n8277, A2 => n8226, ZN => n8275);
   U8363 : NAND2_X1 port map( A1 => n8277, A2 => n8230, ZN => n8278);
   U8364 : NAND2_X1 port map( A1 => n8277, A2 => n8233, ZN => n8280);
   U8365 : NAND2_X1 port map( A1 => n8277, A2 => n8236, ZN => n8282);
   U8366 : NAND2_X1 port map( A1 => n8286, A2 => n8226, ZN => n8284);
   U8367 : NAND2_X1 port map( A1 => n8286, A2 => n8233, ZN => n8289);
   U8368 : NAND2_X1 port map( A1 => n8295, A2 => n8230, ZN => n8296);
   U8369 : NAND2_X1 port map( A1 => n8295, A2 => n8233, ZN => n8298);
   U8370 : NAND2_X1 port map( A1 => n8295, A2 => n8236, ZN => n8300);
   U8371 : NAND2_X1 port map( A1 => n8295, A2 => n8226, ZN => n8293);
   U8372 : NAND2_X1 port map( A1 => n8286, A2 => n8236, ZN => n8291);
   U8373 : NAND2_X1 port map( A1 => n8286, A2 => n8230, ZN => n8287);
   U8374 : NAND2_X1 port map( A1 => n8267, A2 => n8236, ZN => n8272);
   U8375 : NAND2_X1 port map( A1 => n8267, A2 => n8230, ZN => n8268);
   U8376 : NAND2_X1 port map( A1 => n8258, A2 => n8236, ZN => n8263);
   U8377 : NAND2_X1 port map( A1 => n8258, A2 => n8233, ZN => n8261);
   U8378 : NAND2_X1 port map( A1 => n8258, A2 => n8230, ZN => n8259);
   U8379 : NAND2_X1 port map( A1 => n8258, A2 => n8226, ZN => n8256);
   U8380 : NAND2_X1 port map( A1 => n8249, A2 => n8236, ZN => n8254);
   U8381 : NAND2_X1 port map( A1 => n8249, A2 => n8233, ZN => n8252);
   U8382 : NAND2_X1 port map( A1 => n8249, A2 => n8230, ZN => n8250);
   U8383 : NAND2_X1 port map( A1 => n8249, A2 => n8226, ZN => n8247);
   U8384 : NAND2_X1 port map( A1 => n8240, A2 => n8236, ZN => n8245);
   U8385 : NAND2_X1 port map( A1 => n8240, A2 => n8233, ZN => n8243);
   U8386 : NAND2_X1 port map( A1 => n8240, A2 => n8230, ZN => n8241);
   U8387 : NAND2_X1 port map( A1 => n8240, A2 => n8226, ZN => n8238);
   U8388 : NAND2_X1 port map( A1 => n8236, A2 => n8227, ZN => n8234);
   U8389 : NAND2_X1 port map( A1 => n8233, A2 => n8227, ZN => n8231);
   U8390 : NAND2_X1 port map( A1 => n8230, A2 => n8227, ZN => n8228);
   U8391 : NAND2_X1 port map( A1 => n8226, A2 => n8227, ZN => n8224);
   U8392 : AND3_X1 port map( A1 => n8878, A2 => n9686, A3 => n8876, ZN => n8311
                           );
   U8393 : AND3_X1 port map( A1 => n8876, A2 => n9686, A3 => n8877, ZN => n8312
                           );
   U8394 : AND3_X1 port map( A1 => n8875, A2 => n9686, A3 => n8876, ZN => n8316
                           );
   U8395 : AND3_X1 port map( A1 => n8869, A2 => n9687, A3 => n8876, ZN => n8317
                           );
   U8396 : AND3_X1 port map( A1 => n8208, A2 => n10080, A3 => n8209, ZN => 
                           n7644);
   U8397 : AND3_X1 port map( A1 => n8210, A2 => n10080, A3 => n8208, ZN => 
                           n7643);
   U8398 : AND3_X1 port map( A1 => n8201, A2 => n10081, A3 => n8208, ZN => 
                           n7649);
   U8399 : AND3_X1 port map( A1 => n8207, A2 => n10080, A3 => n8208, ZN => 
                           n7648);
   U8400 : AND3_X1 port map( A1 => n8868, A2 => n9686, A3 => n8872, ZN => n8306
                           );
   U8401 : AND3_X1 port map( A1 => n8868, A2 => n9686, A3 => n8871, ZN => n8307
                           );
   U8402 : AND3_X1 port map( A1 => n8200, A2 => n10080, A3 => n8203, ZN => 
                           n7639);
   U8403 : AND3_X1 port map( A1 => n8200, A2 => n10080, A3 => n8204, ZN => 
                           n7638);
   U8404 : AND2_X1 port map( A1 => n8888, A2 => n8877, ZN => n8331);
   U8405 : AND2_X1 port map( A1 => n8887, A2 => n8871, ZN => n8332);
   U8406 : AND2_X1 port map( A1 => n8887, A2 => n8874, ZN => n8342);
   U8407 : AND2_X1 port map( A1 => n8888, A2 => n8874, ZN => n8343);
   U8408 : AND2_X1 port map( A1 => n8888, A2 => n8870, ZN => n8337);
   U8409 : AND2_X1 port map( A1 => n8887, A2 => n8875, ZN => n8338);
   U8410 : AND2_X1 port map( A1 => n8887, A2 => n8872, ZN => n8348);
   U8411 : AND2_X1 port map( A1 => n8888, A2 => n8872, ZN => n8349);
   U8412 : AND2_X1 port map( A1 => n8219, A2 => n8203, ZN => n7664);
   U8413 : AND2_X1 port map( A1 => n8220, A2 => n8209, ZN => n7663);
   U8414 : AND2_X1 port map( A1 => n8220, A2 => n8206, ZN => n7675);
   U8415 : AND2_X1 port map( A1 => n8219, A2 => n8206, ZN => n7674);
   U8416 : AND2_X1 port map( A1 => n8219, A2 => n8207, ZN => n7670);
   U8417 : AND2_X1 port map( A1 => n8220, A2 => n8202, ZN => n7669);
   U8418 : AND2_X1 port map( A1 => n8220, A2 => n8204, ZN => n7681);
   U8419 : AND2_X1 port map( A1 => n8219, A2 => n8204, ZN => n7680);
   U8420 : BUF_X1 port map( A => n6785, Z => n10130);
   U8421 : BUF_X1 port map( A => n6784, Z => n10133);
   U8422 : BUF_X1 port map( A => n6783, Z => n10136);
   U8423 : BUF_X1 port map( A => n6782, Z => n10139);
   U8424 : BUF_X1 port map( A => n6781, Z => n10142);
   U8425 : BUF_X1 port map( A => n6780, Z => n10145);
   U8426 : BUF_X1 port map( A => n6779, Z => n10148);
   U8427 : BUF_X1 port map( A => n6778, Z => n10151);
   U8428 : BUF_X1 port map( A => n6777, Z => n10154);
   U8429 : BUF_X1 port map( A => n6776, Z => n10157);
   U8430 : BUF_X1 port map( A => n6775, Z => n10160);
   U8431 : BUF_X1 port map( A => n6774, Z => n10163);
   U8432 : BUF_X1 port map( A => n6773, Z => n10166);
   U8433 : BUF_X1 port map( A => n6772, Z => n10169);
   U8434 : BUF_X1 port map( A => n6771, Z => n10172);
   U8435 : BUF_X1 port map( A => n6770, Z => n10175);
   U8436 : BUF_X1 port map( A => n6769, Z => n10178);
   U8437 : BUF_X1 port map( A => n6768, Z => n10181);
   U8438 : BUF_X1 port map( A => n6767, Z => n10184);
   U8439 : BUF_X1 port map( A => n6766, Z => n10187);
   U8440 : BUF_X1 port map( A => n6765, Z => n10190);
   U8441 : BUF_X1 port map( A => n6764, Z => n10193);
   U8442 : BUF_X1 port map( A => n6763, Z => n10196);
   U8443 : BUF_X1 port map( A => n6762, Z => n10199);
   U8444 : BUF_X1 port map( A => n6761, Z => n10202);
   U8445 : BUF_X1 port map( A => n6760, Z => n10205);
   U8446 : BUF_X1 port map( A => n6759, Z => n10208);
   U8447 : BUF_X1 port map( A => n6758, Z => n10211);
   U8448 : BUF_X1 port map( A => n6757, Z => n10214);
   U8449 : BUF_X1 port map( A => n6756, Z => n10217);
   U8450 : BUF_X1 port map( A => n6755, Z => n10220);
   U8451 : BUF_X1 port map( A => n6754, Z => n10223);
   U8452 : BUF_X1 port map( A => n6785, Z => n10131);
   U8453 : BUF_X1 port map( A => n6784, Z => n10134);
   U8454 : BUF_X1 port map( A => n6783, Z => n10137);
   U8455 : BUF_X1 port map( A => n6782, Z => n10140);
   U8456 : BUF_X1 port map( A => n6781, Z => n10143);
   U8457 : BUF_X1 port map( A => n6780, Z => n10146);
   U8458 : BUF_X1 port map( A => n6779, Z => n10149);
   U8459 : BUF_X1 port map( A => n6778, Z => n10152);
   U8460 : BUF_X1 port map( A => n6777, Z => n10155);
   U8461 : BUF_X1 port map( A => n6776, Z => n10158);
   U8462 : BUF_X1 port map( A => n6775, Z => n10161);
   U8463 : BUF_X1 port map( A => n6774, Z => n10164);
   U8464 : BUF_X1 port map( A => n6773, Z => n10167);
   U8465 : BUF_X1 port map( A => n6772, Z => n10170);
   U8466 : BUF_X1 port map( A => n6771, Z => n10173);
   U8467 : BUF_X1 port map( A => n6770, Z => n10176);
   U8468 : BUF_X1 port map( A => n6769, Z => n10179);
   U8469 : BUF_X1 port map( A => n6768, Z => n10182);
   U8470 : BUF_X1 port map( A => n6767, Z => n10185);
   U8471 : BUF_X1 port map( A => n6766, Z => n10188);
   U8472 : BUF_X1 port map( A => n6765, Z => n10191);
   U8473 : BUF_X1 port map( A => n6764, Z => n10194);
   U8474 : BUF_X1 port map( A => n6763, Z => n10197);
   U8475 : BUF_X1 port map( A => n6762, Z => n10200);
   U8476 : BUF_X1 port map( A => n6761, Z => n10203);
   U8477 : BUF_X1 port map( A => n6760, Z => n10206);
   U8478 : BUF_X1 port map( A => n6759, Z => n10209);
   U8479 : BUF_X1 port map( A => n6758, Z => n10212);
   U8480 : BUF_X1 port map( A => n6757, Z => n10215);
   U8481 : BUF_X1 port map( A => n6756, Z => n10218);
   U8482 : BUF_X1 port map( A => n6755, Z => n10221);
   U8483 : BUF_X1 port map( A => n6754, Z => n10224);
   U8484 : BUF_X1 port map( A => n9681, Z => n9678);
   U8485 : BUF_X1 port map( A => n9681, Z => n9679);
   U8486 : BUF_X1 port map( A => n10075, Z => n10072);
   U8487 : BUF_X1 port map( A => n10075, Z => n10073);
   U8488 : BUF_X1 port map( A => n6741, Z => n10227);
   U8489 : BUF_X1 port map( A => n6741, Z => n10226);
   U8490 : BUF_X1 port map( A => n9681, Z => n9680);
   U8491 : BUF_X1 port map( A => n10075, Z => n10074);
   U8492 : BUF_X1 port map( A => n6741, Z => n10228);
   U8493 : BUF_X1 port map( A => n6785, Z => n10132);
   U8494 : BUF_X1 port map( A => n6784, Z => n10135);
   U8495 : BUF_X1 port map( A => n6783, Z => n10138);
   U8496 : BUF_X1 port map( A => n6782, Z => n10141);
   U8497 : BUF_X1 port map( A => n6781, Z => n10144);
   U8498 : BUF_X1 port map( A => n6780, Z => n10147);
   U8499 : BUF_X1 port map( A => n6779, Z => n10150);
   U8500 : BUF_X1 port map( A => n6778, Z => n10153);
   U8501 : BUF_X1 port map( A => n6777, Z => n10156);
   U8502 : BUF_X1 port map( A => n6776, Z => n10159);
   U8503 : BUF_X1 port map( A => n6775, Z => n10162);
   U8504 : BUF_X1 port map( A => n6774, Z => n10165);
   U8505 : BUF_X1 port map( A => n6773, Z => n10168);
   U8506 : BUF_X1 port map( A => n6772, Z => n10171);
   U8507 : BUF_X1 port map( A => n6771, Z => n10174);
   U8508 : BUF_X1 port map( A => n6770, Z => n10177);
   U8509 : BUF_X1 port map( A => n6769, Z => n10180);
   U8510 : BUF_X1 port map( A => n6768, Z => n10183);
   U8511 : BUF_X1 port map( A => n6767, Z => n10186);
   U8512 : BUF_X1 port map( A => n6766, Z => n10189);
   U8513 : BUF_X1 port map( A => n6765, Z => n10192);
   U8514 : BUF_X1 port map( A => n6764, Z => n10195);
   U8515 : BUF_X1 port map( A => n6763, Z => n10198);
   U8516 : BUF_X1 port map( A => n6762, Z => n10201);
   U8517 : BUF_X1 port map( A => n6761, Z => n10204);
   U8518 : BUF_X1 port map( A => n6760, Z => n10207);
   U8519 : BUF_X1 port map( A => n6759, Z => n10210);
   U8520 : BUF_X1 port map( A => n6758, Z => n10213);
   U8521 : BUF_X1 port map( A => n6757, Z => n10216);
   U8522 : BUF_X1 port map( A => n6756, Z => n10219);
   U8523 : BUF_X1 port map( A => n6755, Z => n10222);
   U8524 : BUF_X1 port map( A => n6754, Z => n10225);
   U8525 : BUF_X1 port map( A => n9683, Z => n9687);
   U8526 : BUF_X1 port map( A => n9596, Z => n9683);
   U8527 : BUF_X1 port map( A => n10077, Z => n10081);
   U8528 : BUF_X1 port map( A => n9597, Z => n10077);
   U8529 : AOI221_X1 port map( B1 => n9340, B2 => n10061, C1 => n9180, C2 => 
                           n10057, A => n8218, ZN => n8217);
   U8530 : OAI222_X1 port map( A1 => n10053, A2 => n7233, B1 => n10049, B2 => 
                           n6977, C1 => n10045, C2 => n7041, ZN => n8218);
   U8531 : AOI221_X1 port map( B1 => n9341, B2 => n10061, C1 => n9181, C2 => 
                           n10057, A => n8191, ZN => n8190);
   U8532 : OAI222_X1 port map( A1 => n10053, A2 => n7232, B1 => n10049, B2 => 
                           n6976, C1 => n10045, C2 => n7040, ZN => n8191);
   U8533 : AOI221_X1 port map( B1 => n9342, B2 => n10061, C1 => n9182, C2 => 
                           n10057, A => n8174, ZN => n8173);
   U8534 : OAI222_X1 port map( A1 => n10053, A2 => n7231, B1 => n10049, B2 => 
                           n6975, C1 => n10045, C2 => n7039, ZN => n8174);
   U8535 : AOI221_X1 port map( B1 => n9343, B2 => n10061, C1 => n9183, C2 => 
                           n10057, A => n8157, ZN => n8156);
   U8536 : OAI222_X1 port map( A1 => n10053, A2 => n7230, B1 => n10049, B2 => 
                           n6974, C1 => n10045, C2 => n7038, ZN => n8157);
   U8537 : AOI221_X1 port map( B1 => n9344, B2 => n10061, C1 => n9184, C2 => 
                           n10057, A => n8140, ZN => n8139);
   U8538 : OAI222_X1 port map( A1 => n10053, A2 => n7229, B1 => n10049, B2 => 
                           n6973, C1 => n10045, C2 => n7037, ZN => n8140);
   U8539 : AOI221_X1 port map( B1 => n9345, B2 => n10061, C1 => n9185, C2 => 
                           n10057, A => n8123, ZN => n8122);
   U8540 : OAI222_X1 port map( A1 => n10053, A2 => n7228, B1 => n10049, B2 => 
                           n6972, C1 => n10045, C2 => n7036, ZN => n8123);
   U8541 : AOI221_X1 port map( B1 => n9346, B2 => n10061, C1 => n9186, C2 => 
                           n10057, A => n8106, ZN => n8105);
   U8542 : OAI222_X1 port map( A1 => n10053, A2 => n7227, B1 => n10049, B2 => 
                           n6971, C1 => n10045, C2 => n7035, ZN => n8106);
   U8543 : AOI221_X1 port map( B1 => n9347, B2 => n10061, C1 => n9187, C2 => 
                           n10057, A => n8089, ZN => n8088);
   U8544 : OAI222_X1 port map( A1 => n10053, A2 => n7226, B1 => n10049, B2 => 
                           n6970, C1 => n10045, C2 => n7034, ZN => n8089);
   U8545 : AOI221_X1 port map( B1 => n9348, B2 => n10061, C1 => n9188, C2 => 
                           n10057, A => n8072, ZN => n8071);
   U8546 : OAI222_X1 port map( A1 => n10053, A2 => n7225, B1 => n10049, B2 => 
                           n6969, C1 => n10045, C2 => n7033, ZN => n8072);
   U8547 : AOI221_X1 port map( B1 => n9349, B2 => n10061, C1 => n9189, C2 => 
                           n10057, A => n8055, ZN => n8054);
   U8548 : OAI222_X1 port map( A1 => n10053, A2 => n7224, B1 => n10049, B2 => 
                           n6968, C1 => n10045, C2 => n7032, ZN => n8055);
   U8549 : AOI221_X1 port map( B1 => n9350, B2 => n10061, C1 => n9190, C2 => 
                           n10057, A => n8038, ZN => n8037);
   U8550 : OAI222_X1 port map( A1 => n10053, A2 => n7223, B1 => n10049, B2 => 
                           n6967, C1 => n10045, C2 => n7031, ZN => n8038);
   U8551 : AOI221_X1 port map( B1 => n9351, B2 => n10061, C1 => n9191, C2 => 
                           n10057, A => n8021, ZN => n8020);
   U8552 : OAI222_X1 port map( A1 => n10053, A2 => n7222, B1 => n10049, B2 => 
                           n6966, C1 => n10045, C2 => n7030, ZN => n8021);
   U8553 : AOI221_X1 port map( B1 => n9352, B2 => n10062, C1 => n9192, C2 => 
                           n10058, A => n8004, ZN => n8003);
   U8554 : OAI222_X1 port map( A1 => n10054, A2 => n7221, B1 => n10050, B2 => 
                           n6965, C1 => n10046, C2 => n7029, ZN => n8004);
   U8555 : AOI221_X1 port map( B1 => n9353, B2 => n10062, C1 => n9193, C2 => 
                           n10058, A => n7987, ZN => n7986);
   U8556 : OAI222_X1 port map( A1 => n10054, A2 => n7220, B1 => n10050, B2 => 
                           n6964, C1 => n10046, C2 => n7028, ZN => n7987);
   U8557 : AOI221_X1 port map( B1 => n9354, B2 => n10062, C1 => n9194, C2 => 
                           n10058, A => n7970, ZN => n7969);
   U8558 : OAI222_X1 port map( A1 => n10054, A2 => n7219, B1 => n10050, B2 => 
                           n6963, C1 => n10046, C2 => n7027, ZN => n7970);
   U8559 : AOI221_X1 port map( B1 => n9355, B2 => n10062, C1 => n9195, C2 => 
                           n10058, A => n7953, ZN => n7952);
   U8560 : OAI222_X1 port map( A1 => n10054, A2 => n7218, B1 => n10050, B2 => 
                           n6962, C1 => n10046, C2 => n7026, ZN => n7953);
   U8561 : AOI221_X1 port map( B1 => n9356, B2 => n10062, C1 => n9196, C2 => 
                           n10058, A => n7936, ZN => n7935);
   U8562 : OAI222_X1 port map( A1 => n10054, A2 => n7217, B1 => n10050, B2 => 
                           n6961, C1 => n10046, C2 => n7025, ZN => n7936);
   U8563 : AOI221_X1 port map( B1 => n9357, B2 => n10062, C1 => n9197, C2 => 
                           n10058, A => n7919, ZN => n7918);
   U8564 : OAI222_X1 port map( A1 => n10054, A2 => n7216, B1 => n10050, B2 => 
                           n6960, C1 => n10046, C2 => n7024, ZN => n7919);
   U8565 : AOI221_X1 port map( B1 => n9358, B2 => n10062, C1 => n9198, C2 => 
                           n10058, A => n7902, ZN => n7901);
   U8566 : OAI222_X1 port map( A1 => n10054, A2 => n7215, B1 => n10050, B2 => 
                           n6959, C1 => n10046, C2 => n7023, ZN => n7902);
   U8567 : AOI221_X1 port map( B1 => n9359, B2 => n10062, C1 => n9199, C2 => 
                           n10058, A => n7885, ZN => n7884);
   U8568 : OAI222_X1 port map( A1 => n10054, A2 => n7214, B1 => n10050, B2 => 
                           n6958, C1 => n10046, C2 => n7022, ZN => n7885);
   U8569 : AOI221_X1 port map( B1 => n9360, B2 => n10062, C1 => n9200, C2 => 
                           n10058, A => n7868, ZN => n7867);
   U8570 : OAI222_X1 port map( A1 => n10054, A2 => n7213, B1 => n10050, B2 => 
                           n6957, C1 => n10046, C2 => n7021, ZN => n7868);
   U8571 : AOI221_X1 port map( B1 => n9361, B2 => n10062, C1 => n9201, C2 => 
                           n10058, A => n7851, ZN => n7850);
   U8572 : OAI222_X1 port map( A1 => n10054, A2 => n7212, B1 => n10050, B2 => 
                           n6956, C1 => n10046, C2 => n7020, ZN => n7851);
   U8573 : AOI221_X1 port map( B1 => n9362, B2 => n10062, C1 => n9202, C2 => 
                           n10058, A => n7834, ZN => n7833);
   U8574 : OAI222_X1 port map( A1 => n10054, A2 => n7211, B1 => n10050, B2 => 
                           n6955, C1 => n10046, C2 => n7019, ZN => n7834);
   U8575 : AOI221_X1 port map( B1 => n9363, B2 => n10062, C1 => n9203, C2 => 
                           n10058, A => n7817, ZN => n7816);
   U8576 : OAI222_X1 port map( A1 => n10054, A2 => n7210, B1 => n10050, B2 => 
                           n6954, C1 => n10046, C2 => n7018, ZN => n7817);
   U8577 : AOI221_X1 port map( B1 => n9364, B2 => n10063, C1 => n9204, C2 => 
                           n10059, A => n7800, ZN => n7799);
   U8578 : OAI222_X1 port map( A1 => n10055, A2 => n7209, B1 => n10051, B2 => 
                           n6953, C1 => n10047, C2 => n7017, ZN => n7800);
   U8579 : AOI221_X1 port map( B1 => n9365, B2 => n10063, C1 => n9205, C2 => 
                           n10059, A => n7783, ZN => n7782);
   U8580 : OAI222_X1 port map( A1 => n10055, A2 => n7208, B1 => n10051, B2 => 
                           n6952, C1 => n10047, C2 => n7016, ZN => n7783);
   U8581 : AOI221_X1 port map( B1 => n9366, B2 => n10063, C1 => n9206, C2 => 
                           n10059, A => n7766, ZN => n7765);
   U8582 : OAI222_X1 port map( A1 => n10055, A2 => n7207, B1 => n10051, B2 => 
                           n6951, C1 => n10047, C2 => n7015, ZN => n7766);
   U8583 : AOI221_X1 port map( B1 => n9367, B2 => n10063, C1 => n9207, C2 => 
                           n10059, A => n7749, ZN => n7748);
   U8584 : OAI222_X1 port map( A1 => n10055, A2 => n7206, B1 => n10051, B2 => 
                           n6950, C1 => n10047, C2 => n7014, ZN => n7749);
   U8585 : AOI221_X1 port map( B1 => n9368, B2 => n10063, C1 => n9208, C2 => 
                           n10059, A => n7732, ZN => n7731);
   U8586 : OAI222_X1 port map( A1 => n10055, A2 => n7205, B1 => n10051, B2 => 
                           n6949, C1 => n10047, C2 => n7013, ZN => n7732);
   U8587 : AOI221_X1 port map( B1 => n9369, B2 => n10063, C1 => n9209, C2 => 
                           n10059, A => n7715, ZN => n7714);
   U8588 : OAI222_X1 port map( A1 => n10055, A2 => n7204, B1 => n10051, B2 => 
                           n6948, C1 => n10047, C2 => n7012, ZN => n7715);
   U8589 : AOI221_X1 port map( B1 => n9370, B2 => n10063, C1 => n9210, C2 => 
                           n10059, A => n7698, ZN => n7697);
   U8590 : OAI222_X1 port map( A1 => n10055, A2 => n7203, B1 => n10051, B2 => 
                           n6947, C1 => n10047, C2 => n7011, ZN => n7698);
   U8591 : AOI221_X1 port map( B1 => n9371, B2 => n10063, C1 => n9211, C2 => 
                           n10059, A => n7665, ZN => n7662);
   U8592 : OAI222_X1 port map( A1 => n10055, A2 => n7202, B1 => n10051, B2 => 
                           n6946, C1 => n10047, C2 => n7010, ZN => n7665);
   U8593 : AOI221_X1 port map( B1 => n10078, B2 => n8212, C1 => n10072, C2 => 
                           OUT2_0_port, A => n8213, ZN => n8195);
   U8594 : OAI22_X1 port map( A1 => n10068, A2 => n7456, B1 => n10064, B2 => 
                           n7424, ZN => n8213);
   U8595 : NAND4_X1 port map( A1 => n8214, A2 => n8215, A3 => n8216, A4 => 
                           n8217, ZN => n8212);
   U8596 : AOI221_X1 port map( B1 => n9148, B2 => n10005, C1 => n9020, C2 => 
                           n10001, A => n8223, ZN => n8214);
   U8597 : AOI221_X1 port map( B1 => n10080, B2 => n8185, C1 => n10072, C2 => 
                           OUT2_1_port, A => n8186, ZN => n8178);
   U8598 : OAI22_X1 port map( A1 => n10068, A2 => n7455, B1 => n10064, B2 => 
                           n7423, ZN => n8186);
   U8599 : NAND4_X1 port map( A1 => n8187, A2 => n8188, A3 => n8189, A4 => 
                           n8190, ZN => n8185);
   U8600 : AOI221_X1 port map( B1 => n9149, B2 => n10005, C1 => n9021, C2 => 
                           n10001, A => n8194, ZN => n8187);
   U8601 : AOI221_X1 port map( B1 => n10080, B2 => n8168, C1 => n10072, C2 => 
                           OUT2_2_port, A => n8169, ZN => n8161);
   U8602 : OAI22_X1 port map( A1 => n10068, A2 => n7454, B1 => n10064, B2 => 
                           n7422, ZN => n8169);
   U8603 : NAND4_X1 port map( A1 => n8170, A2 => n8171, A3 => n8172, A4 => 
                           n8173, ZN => n8168);
   U8604 : AOI221_X1 port map( B1 => n9150, B2 => n10005, C1 => n9022, C2 => 
                           n10001, A => n8177, ZN => n8170);
   U8605 : AOI221_X1 port map( B1 => n10079, B2 => n8151, C1 => n10072, C2 => 
                           OUT2_3_port, A => n8152, ZN => n8144);
   U8606 : OAI22_X1 port map( A1 => n10068, A2 => n7453, B1 => n10064, B2 => 
                           n7421, ZN => n8152);
   U8607 : NAND4_X1 port map( A1 => n8153, A2 => n8154, A3 => n8155, A4 => 
                           n8156, ZN => n8151);
   U8608 : AOI221_X1 port map( B1 => n9151, B2 => n10005, C1 => n9023, C2 => 
                           n10001, A => n8160, ZN => n8153);
   U8609 : AOI221_X1 port map( B1 => n10080, B2 => n8134, C1 => n10072, C2 => 
                           OUT2_4_port, A => n8135, ZN => n8127);
   U8610 : OAI22_X1 port map( A1 => n10068, A2 => n7452, B1 => n10064, B2 => 
                           n7420, ZN => n8135);
   U8611 : NAND4_X1 port map( A1 => n8136, A2 => n8137, A3 => n8138, A4 => 
                           n8139, ZN => n8134);
   U8612 : AOI221_X1 port map( B1 => n9152, B2 => n10005, C1 => n9024, C2 => 
                           n10001, A => n8143, ZN => n8136);
   U8613 : AOI221_X1 port map( B1 => n10080, B2 => n8117, C1 => n10072, C2 => 
                           OUT2_5_port, A => n8118, ZN => n8110);
   U8614 : OAI22_X1 port map( A1 => n10068, A2 => n7451, B1 => n10064, B2 => 
                           n7419, ZN => n8118);
   U8615 : NAND4_X1 port map( A1 => n8119, A2 => n8120, A3 => n8121, A4 => 
                           n8122, ZN => n8117);
   U8616 : AOI221_X1 port map( B1 => n9153, B2 => n10005, C1 => n9025, C2 => 
                           n10001, A => n8126, ZN => n8119);
   U8617 : AOI221_X1 port map( B1 => n10080, B2 => n8100, C1 => n10072, C2 => 
                           OUT2_6_port, A => n8101, ZN => n8093);
   U8618 : OAI22_X1 port map( A1 => n10068, A2 => n7450, B1 => n10064, B2 => 
                           n7418, ZN => n8101);
   U8619 : NAND4_X1 port map( A1 => n8102, A2 => n8103, A3 => n8104, A4 => 
                           n8105, ZN => n8100);
   U8620 : AOI221_X1 port map( B1 => n9154, B2 => n10005, C1 => n9026, C2 => 
                           n10001, A => n8109, ZN => n8102);
   U8621 : AOI221_X1 port map( B1 => n10080, B2 => n8083, C1 => n10072, C2 => 
                           OUT2_7_port, A => n8084, ZN => n8076);
   U8622 : OAI22_X1 port map( A1 => n10068, A2 => n7449, B1 => n10064, B2 => 
                           n7417, ZN => n8084);
   U8623 : NAND4_X1 port map( A1 => n8085, A2 => n8086, A3 => n8087, A4 => 
                           n8088, ZN => n8083);
   U8624 : AOI221_X1 port map( B1 => n9155, B2 => n10005, C1 => n9027, C2 => 
                           n10001, A => n8092, ZN => n8085);
   U8625 : AOI221_X1 port map( B1 => n10080, B2 => n8066, C1 => n10072, C2 => 
                           OUT2_8_port, A => n8067, ZN => n8059);
   U8626 : OAI22_X1 port map( A1 => n10068, A2 => n7448, B1 => n10064, B2 => 
                           n7416, ZN => n8067);
   U8627 : NAND4_X1 port map( A1 => n8068, A2 => n8069, A3 => n8070, A4 => 
                           n8071, ZN => n8066);
   U8628 : AOI221_X1 port map( B1 => n9156, B2 => n10005, C1 => n9028, C2 => 
                           n10001, A => n8075, ZN => n8068);
   U8629 : AOI221_X1 port map( B1 => n10080, B2 => n8049, C1 => n10072, C2 => 
                           OUT2_9_port, A => n8050, ZN => n8042);
   U8630 : OAI22_X1 port map( A1 => n10068, A2 => n7447, B1 => n10064, B2 => 
                           n7415, ZN => n8050);
   U8631 : NAND4_X1 port map( A1 => n8051, A2 => n8052, A3 => n8053, A4 => 
                           n8054, ZN => n8049);
   U8632 : AOI221_X1 port map( B1 => n9157, B2 => n10005, C1 => n9029, C2 => 
                           n10001, A => n8058, ZN => n8051);
   U8633 : AOI221_X1 port map( B1 => n10080, B2 => n8032, C1 => n10072, C2 => 
                           OUT2_10_port, A => n8033, ZN => n8025);
   U8634 : OAI22_X1 port map( A1 => n10068, A2 => n7446, B1 => n10064, B2 => 
                           n7414, ZN => n8033);
   U8635 : NAND4_X1 port map( A1 => n8034, A2 => n8035, A3 => n8036, A4 => 
                           n8037, ZN => n8032);
   U8636 : AOI221_X1 port map( B1 => n9158, B2 => n10005, C1 => n9030, C2 => 
                           n10001, A => n8041, ZN => n8034);
   U8637 : AOI221_X1 port map( B1 => n10079, B2 => n8015, C1 => n10072, C2 => 
                           OUT2_11_port, A => n8016, ZN => n8008);
   U8638 : OAI22_X1 port map( A1 => n10068, A2 => n7445, B1 => n10064, B2 => 
                           n7413, ZN => n8016);
   U8639 : NAND4_X1 port map( A1 => n8017, A2 => n8018, A3 => n8019, A4 => 
                           n8020, ZN => n8015);
   U8640 : AOI221_X1 port map( B1 => n9159, B2 => n10005, C1 => n9031, C2 => 
                           n10001, A => n8024, ZN => n8017);
   U8641 : AOI221_X1 port map( B1 => n10079, B2 => n7998, C1 => n10073, C2 => 
                           OUT2_12_port, A => n7999, ZN => n7991);
   U8642 : OAI22_X1 port map( A1 => n10069, A2 => n7444, B1 => n10065, B2 => 
                           n7412, ZN => n7999);
   U8643 : NAND4_X1 port map( A1 => n8000, A2 => n8001, A3 => n8002, A4 => 
                           n8003, ZN => n7998);
   U8644 : AOI221_X1 port map( B1 => n9160, B2 => n10006, C1 => n9032, C2 => 
                           n10002, A => n8007, ZN => n8000);
   U8645 : AOI221_X1 port map( B1 => n10079, B2 => n7981, C1 => n10073, C2 => 
                           OUT2_13_port, A => n7982, ZN => n7974);
   U8646 : OAI22_X1 port map( A1 => n10069, A2 => n7443, B1 => n10065, B2 => 
                           n7411, ZN => n7982);
   U8647 : NAND4_X1 port map( A1 => n7983, A2 => n7984, A3 => n7985, A4 => 
                           n7986, ZN => n7981);
   U8648 : AOI221_X1 port map( B1 => n9161, B2 => n10006, C1 => n9033, C2 => 
                           n10002, A => n7990, ZN => n7983);
   U8649 : AOI221_X1 port map( B1 => n10079, B2 => n7964, C1 => n10073, C2 => 
                           OUT2_14_port, A => n7965, ZN => n7957);
   U8650 : OAI22_X1 port map( A1 => n10069, A2 => n7442, B1 => n10065, B2 => 
                           n7410, ZN => n7965);
   U8651 : NAND4_X1 port map( A1 => n7966, A2 => n7967, A3 => n7968, A4 => 
                           n7969, ZN => n7964);
   U8652 : AOI221_X1 port map( B1 => n9162, B2 => n10006, C1 => n9034, C2 => 
                           n10002, A => n7973, ZN => n7966);
   U8653 : AOI221_X1 port map( B1 => n10079, B2 => n7947, C1 => n10073, C2 => 
                           OUT2_15_port, A => n7948, ZN => n7940);
   U8654 : OAI22_X1 port map( A1 => n10069, A2 => n7441, B1 => n10065, B2 => 
                           n7409, ZN => n7948);
   U8655 : NAND4_X1 port map( A1 => n7949, A2 => n7950, A3 => n7951, A4 => 
                           n7952, ZN => n7947);
   U8656 : AOI221_X1 port map( B1 => n9163, B2 => n10006, C1 => n9035, C2 => 
                           n10002, A => n7956, ZN => n7949);
   U8657 : AOI221_X1 port map( B1 => n10079, B2 => n7930, C1 => n10073, C2 => 
                           OUT2_16_port, A => n7931, ZN => n7923);
   U8658 : OAI22_X1 port map( A1 => n10069, A2 => n7440, B1 => n10065, B2 => 
                           n7408, ZN => n7931);
   U8659 : NAND4_X1 port map( A1 => n7932, A2 => n7933, A3 => n7934, A4 => 
                           n7935, ZN => n7930);
   U8660 : AOI221_X1 port map( B1 => n9164, B2 => n10006, C1 => n9036, C2 => 
                           n10002, A => n7939, ZN => n7932);
   U8661 : AOI221_X1 port map( B1 => n10079, B2 => n7913, C1 => n10073, C2 => 
                           OUT2_17_port, A => n7914, ZN => n7906);
   U8662 : OAI22_X1 port map( A1 => n10069, A2 => n7439, B1 => n10065, B2 => 
                           n7407, ZN => n7914);
   U8663 : NAND4_X1 port map( A1 => n7915, A2 => n7916, A3 => n7917, A4 => 
                           n7918, ZN => n7913);
   U8664 : AOI221_X1 port map( B1 => n9165, B2 => n10006, C1 => n9037, C2 => 
                           n10002, A => n7922, ZN => n7915);
   U8665 : AOI221_X1 port map( B1 => n10079, B2 => n7896, C1 => n10073, C2 => 
                           OUT2_18_port, A => n7897, ZN => n7889);
   U8666 : OAI22_X1 port map( A1 => n10069, A2 => n7438, B1 => n10065, B2 => 
                           n7406, ZN => n7897);
   U8667 : NAND4_X1 port map( A1 => n7898, A2 => n7899, A3 => n7900, A4 => 
                           n7901, ZN => n7896);
   U8668 : AOI221_X1 port map( B1 => n9166, B2 => n10006, C1 => n9038, C2 => 
                           n10002, A => n7905, ZN => n7898);
   U8669 : AOI221_X1 port map( B1 => n10079, B2 => n7879, C1 => n10073, C2 => 
                           OUT2_19_port, A => n7880, ZN => n7872);
   U8670 : OAI22_X1 port map( A1 => n10069, A2 => n7437, B1 => n10065, B2 => 
                           n7405, ZN => n7880);
   U8671 : NAND4_X1 port map( A1 => n7881, A2 => n7882, A3 => n7883, A4 => 
                           n7884, ZN => n7879);
   U8672 : AOI221_X1 port map( B1 => n9167, B2 => n10006, C1 => n9039, C2 => 
                           n10002, A => n7888, ZN => n7881);
   U8673 : AOI221_X1 port map( B1 => n10079, B2 => n7862, C1 => n10073, C2 => 
                           OUT2_20_port, A => n7863, ZN => n7855);
   U8674 : OAI22_X1 port map( A1 => n10069, A2 => n7436, B1 => n10065, B2 => 
                           n7404, ZN => n7863);
   U8675 : NAND4_X1 port map( A1 => n7864, A2 => n7865, A3 => n7866, A4 => 
                           n7867, ZN => n7862);
   U8676 : AOI221_X1 port map( B1 => n9168, B2 => n10006, C1 => n9040, C2 => 
                           n10002, A => n7871, ZN => n7864);
   U8677 : AOI221_X1 port map( B1 => n10079, B2 => n7845, C1 => n10073, C2 => 
                           OUT2_21_port, A => n7846, ZN => n7838);
   U8678 : OAI22_X1 port map( A1 => n10069, A2 => n7435, B1 => n10065, B2 => 
                           n7403, ZN => n7846);
   U8679 : NAND4_X1 port map( A1 => n7847, A2 => n7848, A3 => n7849, A4 => 
                           n7850, ZN => n7845);
   U8680 : AOI221_X1 port map( B1 => n9169, B2 => n10006, C1 => n9041, C2 => 
                           n10002, A => n7854, ZN => n7847);
   U8681 : AOI221_X1 port map( B1 => n10078, B2 => n7828, C1 => n10073, C2 => 
                           OUT2_22_port, A => n7829, ZN => n7821);
   U8682 : OAI22_X1 port map( A1 => n10069, A2 => n7434, B1 => n10065, B2 => 
                           n7402, ZN => n7829);
   U8683 : NAND4_X1 port map( A1 => n7830, A2 => n7831, A3 => n7832, A4 => 
                           n7833, ZN => n7828);
   U8684 : AOI221_X1 port map( B1 => n9170, B2 => n10006, C1 => n9042, C2 => 
                           n10002, A => n7837, ZN => n7830);
   U8685 : AOI221_X1 port map( B1 => n10078, B2 => n7811, C1 => n10073, C2 => 
                           OUT2_23_port, A => n7812, ZN => n7804);
   U8686 : OAI22_X1 port map( A1 => n10069, A2 => n7433, B1 => n10065, B2 => 
                           n7401, ZN => n7812);
   U8687 : NAND4_X1 port map( A1 => n7813, A2 => n7814, A3 => n7815, A4 => 
                           n7816, ZN => n7811);
   U8688 : AOI221_X1 port map( B1 => n9171, B2 => n10006, C1 => n9043, C2 => 
                           n10002, A => n7820, ZN => n7813);
   U8689 : AOI221_X1 port map( B1 => n10078, B2 => n7794, C1 => n10074, C2 => 
                           OUT2_24_port, A => n7795, ZN => n7787);
   U8690 : OAI22_X1 port map( A1 => n10070, A2 => n7432, B1 => n10066, B2 => 
                           n7400, ZN => n7795);
   U8691 : NAND4_X1 port map( A1 => n7796, A2 => n7797, A3 => n7798, A4 => 
                           n7799, ZN => n7794);
   U8692 : AOI221_X1 port map( B1 => n9172, B2 => n10007, C1 => n9044, C2 => 
                           n10003, A => n7803, ZN => n7796);
   U8693 : AOI221_X1 port map( B1 => n10078, B2 => n7777, C1 => n10074, C2 => 
                           OUT2_25_port, A => n7778, ZN => n7770);
   U8694 : OAI22_X1 port map( A1 => n10070, A2 => n7431, B1 => n10066, B2 => 
                           n7399, ZN => n7778);
   U8695 : NAND4_X1 port map( A1 => n7779, A2 => n7780, A3 => n7781, A4 => 
                           n7782, ZN => n7777);
   U8696 : AOI221_X1 port map( B1 => n9173, B2 => n10007, C1 => n9045, C2 => 
                           n10003, A => n7786, ZN => n7779);
   U8697 : AOI221_X1 port map( B1 => n10078, B2 => n7760, C1 => n10074, C2 => 
                           OUT2_26_port, A => n7761, ZN => n7753);
   U8698 : OAI22_X1 port map( A1 => n10070, A2 => n7430, B1 => n10066, B2 => 
                           n7398, ZN => n7761);
   U8699 : NAND4_X1 port map( A1 => n7762, A2 => n7763, A3 => n7764, A4 => 
                           n7765, ZN => n7760);
   U8700 : AOI221_X1 port map( B1 => n9174, B2 => n10007, C1 => n9046, C2 => 
                           n10003, A => n7769, ZN => n7762);
   U8701 : AOI221_X1 port map( B1 => n10078, B2 => n7743, C1 => n10074, C2 => 
                           OUT2_27_port, A => n7744, ZN => n7736);
   U8702 : OAI22_X1 port map( A1 => n10070, A2 => n7429, B1 => n10066, B2 => 
                           n7397, ZN => n7744);
   U8703 : NAND4_X1 port map( A1 => n7745, A2 => n7746, A3 => n7747, A4 => 
                           n7748, ZN => n7743);
   U8704 : AOI221_X1 port map( B1 => n9175, B2 => n10007, C1 => n9047, C2 => 
                           n10003, A => n7752, ZN => n7745);
   U8705 : AOI221_X1 port map( B1 => n10078, B2 => n7726, C1 => n10074, C2 => 
                           OUT2_28_port, A => n7727, ZN => n7719);
   U8706 : OAI22_X1 port map( A1 => n10070, A2 => n7428, B1 => n10066, B2 => 
                           n7396, ZN => n7727);
   U8707 : NAND4_X1 port map( A1 => n7728, A2 => n7729, A3 => n7730, A4 => 
                           n7731, ZN => n7726);
   U8708 : AOI221_X1 port map( B1 => n9176, B2 => n10007, C1 => n9048, C2 => 
                           n10003, A => n7735, ZN => n7728);
   U8709 : AOI221_X1 port map( B1 => n10078, B2 => n7709, C1 => n10074, C2 => 
                           OUT2_29_port, A => n7710, ZN => n7702);
   U8710 : OAI22_X1 port map( A1 => n10070, A2 => n7427, B1 => n10066, B2 => 
                           n7395, ZN => n7710);
   U8711 : NAND4_X1 port map( A1 => n7711, A2 => n7712, A3 => n7713, A4 => 
                           n7714, ZN => n7709);
   U8712 : AOI221_X1 port map( B1 => n9177, B2 => n10007, C1 => n9049, C2 => 
                           n10003, A => n7718, ZN => n7711);
   U8713 : AOI221_X1 port map( B1 => n10078, B2 => n7692, C1 => n10074, C2 => 
                           OUT2_30_port, A => n7693, ZN => n7685);
   U8714 : OAI22_X1 port map( A1 => n10070, A2 => n7426, B1 => n10066, B2 => 
                           n7394, ZN => n7693);
   U8715 : NAND4_X1 port map( A1 => n7694, A2 => n7695, A3 => n7696, A4 => 
                           n7697, ZN => n7692);
   U8716 : AOI221_X1 port map( B1 => n9178, B2 => n10007, C1 => n9050, C2 => 
                           n10003, A => n7701, ZN => n7694);
   U8717 : AOI221_X1 port map( B1 => n10078, B2 => n7654, C1 => n10074, C2 => 
                           OUT2_31_port, A => n7656, ZN => n7634);
   U8718 : OAI22_X1 port map( A1 => n10070, A2 => n7425, B1 => n10066, B2 => 
                           n7393, ZN => n7656);
   U8719 : NAND4_X1 port map( A1 => n7659, A2 => n7660, A3 => n7661, A4 => 
                           n7662, ZN => n7654);
   U8720 : AOI221_X1 port map( B1 => n9179, B2 => n10007, C1 => n9051, C2 => 
                           n10003, A => n7682, ZN => n7659);
   U8721 : NAND4_X1 port map( A1 => n8195, A2 => n8196, A3 => n8197, A4 => 
                           n8198, ZN => n2336);
   U8722 : AOI221_X1 port map( B1 => n10127, B2 => n7632, C1 => n9308, C2 => 
                           n10123, A => n8199, ZN => n8198);
   U8723 : AOI221_X1 port map( B1 => n4679, B2 => n10095, C1 => n4743, C2 => 
                           n10091, A => n8211, ZN => n8196);
   U8724 : AOI221_X1 port map( B1 => n4711, B2 => n10111, C1 => n9244, C2 => 
                           n10107, A => n8205, ZN => n8197);
   U8725 : NAND4_X1 port map( A1 => n8178, A2 => n8179, A3 => n8180, A4 => 
                           n8181, ZN => n2337);
   U8726 : AOI221_X1 port map( B1 => n10127, B2 => n7631, C1 => n9309, C2 => 
                           n10123, A => n8182, ZN => n8181);
   U8727 : AOI221_X1 port map( B1 => n4678, B2 => n10095, C1 => n4742, C2 => 
                           n10091, A => n8184, ZN => n8179);
   U8728 : AOI221_X1 port map( B1 => n4710, B2 => n10111, C1 => n9245, C2 => 
                           n10107, A => n8183, ZN => n8180);
   U8729 : NAND4_X1 port map( A1 => n8161, A2 => n8162, A3 => n8163, A4 => 
                           n8164, ZN => n2338);
   U8730 : AOI221_X1 port map( B1 => n10127, B2 => n7630, C1 => n9310, C2 => 
                           n10123, A => n8165, ZN => n8164);
   U8731 : AOI221_X1 port map( B1 => n4677, B2 => n10095, C1 => n4741, C2 => 
                           n10091, A => n8167, ZN => n8162);
   U8732 : AOI221_X1 port map( B1 => n4709, B2 => n10111, C1 => n9246, C2 => 
                           n10107, A => n8166, ZN => n8163);
   U8733 : NAND4_X1 port map( A1 => n8144, A2 => n8145, A3 => n8146, A4 => 
                           n8147, ZN => n2339);
   U8734 : AOI221_X1 port map( B1 => n10127, B2 => n7629, C1 => n9311, C2 => 
                           n10123, A => n8148, ZN => n8147);
   U8735 : AOI221_X1 port map( B1 => n4676, B2 => n10095, C1 => n4740, C2 => 
                           n10091, A => n8150, ZN => n8145);
   U8736 : AOI221_X1 port map( B1 => n4708, B2 => n10111, C1 => n9247, C2 => 
                           n10107, A => n8149, ZN => n8146);
   U8737 : NAND4_X1 port map( A1 => n8127, A2 => n8128, A3 => n8129, A4 => 
                           n8130, ZN => n2340);
   U8738 : AOI221_X1 port map( B1 => n10127, B2 => n7628, C1 => n9312, C2 => 
                           n10123, A => n8131, ZN => n8130);
   U8739 : AOI221_X1 port map( B1 => n4675, B2 => n10095, C1 => n4739, C2 => 
                           n10091, A => n8133, ZN => n8128);
   U8740 : AOI221_X1 port map( B1 => n4707, B2 => n10111, C1 => n9248, C2 => 
                           n10107, A => n8132, ZN => n8129);
   U8741 : NAND4_X1 port map( A1 => n8110, A2 => n8111, A3 => n8112, A4 => 
                           n8113, ZN => n2341);
   U8742 : AOI221_X1 port map( B1 => n10127, B2 => n7627, C1 => n9313, C2 => 
                           n10123, A => n8114, ZN => n8113);
   U8743 : AOI221_X1 port map( B1 => n4674, B2 => n10095, C1 => n4738, C2 => 
                           n10091, A => n8116, ZN => n8111);
   U8744 : AOI221_X1 port map( B1 => n4706, B2 => n10111, C1 => n9249, C2 => 
                           n10107, A => n8115, ZN => n8112);
   U8745 : NAND4_X1 port map( A1 => n8093, A2 => n8094, A3 => n8095, A4 => 
                           n8096, ZN => n2342);
   U8746 : AOI221_X1 port map( B1 => n10127, B2 => n7626, C1 => n9314, C2 => 
                           n10123, A => n8097, ZN => n8096);
   U8747 : AOI221_X1 port map( B1 => n4673, B2 => n10095, C1 => n4737, C2 => 
                           n10091, A => n8099, ZN => n8094);
   U8748 : AOI221_X1 port map( B1 => n4705, B2 => n10111, C1 => n9250, C2 => 
                           n10107, A => n8098, ZN => n8095);
   U8749 : NAND4_X1 port map( A1 => n8076, A2 => n8077, A3 => n8078, A4 => 
                           n8079, ZN => n2343);
   U8750 : AOI221_X1 port map( B1 => n10127, B2 => n7625, C1 => n9315, C2 => 
                           n10123, A => n8080, ZN => n8079);
   U8751 : AOI221_X1 port map( B1 => n4672, B2 => n10095, C1 => n4736, C2 => 
                           n10091, A => n8082, ZN => n8077);
   U8752 : AOI221_X1 port map( B1 => n4704, B2 => n10111, C1 => n9251, C2 => 
                           n10107, A => n8081, ZN => n8078);
   U8753 : NAND4_X1 port map( A1 => n8059, A2 => n8060, A3 => n8061, A4 => 
                           n8062, ZN => n2344);
   U8754 : AOI221_X1 port map( B1 => n10127, B2 => n7624, C1 => n9316, C2 => 
                           n10123, A => n8063, ZN => n8062);
   U8755 : AOI221_X1 port map( B1 => n4671, B2 => n10095, C1 => n4735, C2 => 
                           n10091, A => n8065, ZN => n8060);
   U8756 : AOI221_X1 port map( B1 => n4703, B2 => n10111, C1 => n9252, C2 => 
                           n10107, A => n8064, ZN => n8061);
   U8757 : NAND4_X1 port map( A1 => n8042, A2 => n8043, A3 => n8044, A4 => 
                           n8045, ZN => n2345);
   U8758 : AOI221_X1 port map( B1 => n10127, B2 => n7623, C1 => n9317, C2 => 
                           n10123, A => n8046, ZN => n8045);
   U8759 : AOI221_X1 port map( B1 => n4670, B2 => n10095, C1 => n4734, C2 => 
                           n10091, A => n8048, ZN => n8043);
   U8760 : AOI221_X1 port map( B1 => n4702, B2 => n10111, C1 => n9253, C2 => 
                           n10107, A => n8047, ZN => n8044);
   U8761 : NAND4_X1 port map( A1 => n8025, A2 => n8026, A3 => n8027, A4 => 
                           n8028, ZN => n2346);
   U8762 : AOI221_X1 port map( B1 => n10127, B2 => n7622, C1 => n9318, C2 => 
                           n10123, A => n8029, ZN => n8028);
   U8763 : AOI221_X1 port map( B1 => n4669, B2 => n10095, C1 => n4733, C2 => 
                           n10091, A => n8031, ZN => n8026);
   U8764 : AOI221_X1 port map( B1 => n4701, B2 => n10111, C1 => n9254, C2 => 
                           n10107, A => n8030, ZN => n8027);
   U8765 : NAND4_X1 port map( A1 => n8008, A2 => n8009, A3 => n8010, A4 => 
                           n8011, ZN => n2347);
   U8766 : AOI221_X1 port map( B1 => n10127, B2 => n7621, C1 => n9319, C2 => 
                           n10123, A => n8012, ZN => n8011);
   U8767 : AOI221_X1 port map( B1 => n4668, B2 => n10095, C1 => n4732, C2 => 
                           n10091, A => n8014, ZN => n8009);
   U8768 : AOI221_X1 port map( B1 => n4700, B2 => n10111, C1 => n9255, C2 => 
                           n10107, A => n8013, ZN => n8010);
   U8769 : NAND4_X1 port map( A1 => n7991, A2 => n7992, A3 => n7993, A4 => 
                           n7994, ZN => n2348);
   U8770 : AOI221_X1 port map( B1 => n10128, B2 => n7620, C1 => n9320, C2 => 
                           n10124, A => n7995, ZN => n7994);
   U8771 : AOI221_X1 port map( B1 => n4667, B2 => n10096, C1 => n4731, C2 => 
                           n10092, A => n7997, ZN => n7992);
   U8772 : AOI221_X1 port map( B1 => n4699, B2 => n10112, C1 => n9256, C2 => 
                           n10108, A => n7996, ZN => n7993);
   U8773 : NAND4_X1 port map( A1 => n7974, A2 => n7975, A3 => n7976, A4 => 
                           n7977, ZN => n2349);
   U8774 : AOI221_X1 port map( B1 => n10128, B2 => n7619, C1 => n9321, C2 => 
                           n10124, A => n7978, ZN => n7977);
   U8775 : AOI221_X1 port map( B1 => n4666, B2 => n10096, C1 => n4730, C2 => 
                           n10092, A => n7980, ZN => n7975);
   U8776 : AOI221_X1 port map( B1 => n4698, B2 => n10112, C1 => n9257, C2 => 
                           n10108, A => n7979, ZN => n7976);
   U8777 : NAND4_X1 port map( A1 => n7957, A2 => n7958, A3 => n7959, A4 => 
                           n7960, ZN => n2350);
   U8778 : AOI221_X1 port map( B1 => n10128, B2 => n7618, C1 => n9322, C2 => 
                           n10124, A => n7961, ZN => n7960);
   U8779 : AOI221_X1 port map( B1 => n4665, B2 => n10096, C1 => n4729, C2 => 
                           n10092, A => n7963, ZN => n7958);
   U8780 : AOI221_X1 port map( B1 => n4697, B2 => n10112, C1 => n9258, C2 => 
                           n10108, A => n7962, ZN => n7959);
   U8781 : NAND4_X1 port map( A1 => n7940, A2 => n7941, A3 => n7942, A4 => 
                           n7943, ZN => n2351);
   U8782 : AOI221_X1 port map( B1 => n10128, B2 => n7617, C1 => n9323, C2 => 
                           n10124, A => n7944, ZN => n7943);
   U8783 : AOI221_X1 port map( B1 => n4664, B2 => n10096, C1 => n4728, C2 => 
                           n10092, A => n7946, ZN => n7941);
   U8784 : AOI221_X1 port map( B1 => n4696, B2 => n10112, C1 => n9259, C2 => 
                           n10108, A => n7945, ZN => n7942);
   U8785 : NAND4_X1 port map( A1 => n7923, A2 => n7924, A3 => n7925, A4 => 
                           n7926, ZN => n2352);
   U8786 : AOI221_X1 port map( B1 => n10128, B2 => n7616, C1 => n9324, C2 => 
                           n10124, A => n7927, ZN => n7926);
   U8787 : AOI221_X1 port map( B1 => n4663, B2 => n10096, C1 => n4727, C2 => 
                           n10092, A => n7929, ZN => n7924);
   U8788 : AOI221_X1 port map( B1 => n4695, B2 => n10112, C1 => n9260, C2 => 
                           n10108, A => n7928, ZN => n7925);
   U8789 : NAND4_X1 port map( A1 => n7906, A2 => n7907, A3 => n7908, A4 => 
                           n7909, ZN => n2353);
   U8790 : AOI221_X1 port map( B1 => n10128, B2 => n7615, C1 => n9325, C2 => 
                           n10124, A => n7910, ZN => n7909);
   U8791 : AOI221_X1 port map( B1 => n4662, B2 => n10096, C1 => n4726, C2 => 
                           n10092, A => n7912, ZN => n7907);
   U8792 : AOI221_X1 port map( B1 => n4694, B2 => n10112, C1 => n9261, C2 => 
                           n10108, A => n7911, ZN => n7908);
   U8793 : NAND4_X1 port map( A1 => n7889, A2 => n7890, A3 => n7891, A4 => 
                           n7892, ZN => n2354);
   U8794 : AOI221_X1 port map( B1 => n10128, B2 => n7614, C1 => n9326, C2 => 
                           n10124, A => n7893, ZN => n7892);
   U8795 : AOI221_X1 port map( B1 => n4661, B2 => n10096, C1 => n4725, C2 => 
                           n10092, A => n7895, ZN => n7890);
   U8796 : AOI221_X1 port map( B1 => n4693, B2 => n10112, C1 => n9262, C2 => 
                           n10108, A => n7894, ZN => n7891);
   U8797 : NAND4_X1 port map( A1 => n7872, A2 => n7873, A3 => n7874, A4 => 
                           n7875, ZN => n2355);
   U8798 : AOI221_X1 port map( B1 => n10128, B2 => n7613, C1 => n9327, C2 => 
                           n10124, A => n7876, ZN => n7875);
   U8799 : AOI221_X1 port map( B1 => n4660, B2 => n10096, C1 => n4724, C2 => 
                           n10092, A => n7878, ZN => n7873);
   U8800 : AOI221_X1 port map( B1 => n4692, B2 => n10112, C1 => n9263, C2 => 
                           n10108, A => n7877, ZN => n7874);
   U8801 : NAND4_X1 port map( A1 => n7855, A2 => n7856, A3 => n7857, A4 => 
                           n7858, ZN => n2356);
   U8802 : AOI221_X1 port map( B1 => n10128, B2 => n7612, C1 => n9328, C2 => 
                           n10124, A => n7859, ZN => n7858);
   U8803 : AOI221_X1 port map( B1 => n4659, B2 => n10096, C1 => n4723, C2 => 
                           n10092, A => n7861, ZN => n7856);
   U8804 : AOI221_X1 port map( B1 => n4691, B2 => n10112, C1 => n9264, C2 => 
                           n10108, A => n7860, ZN => n7857);
   U8805 : NAND4_X1 port map( A1 => n7838, A2 => n7839, A3 => n7840, A4 => 
                           n7841, ZN => n2357);
   U8806 : AOI221_X1 port map( B1 => n10128, B2 => n7611, C1 => n9329, C2 => 
                           n10124, A => n7842, ZN => n7841);
   U8807 : AOI221_X1 port map( B1 => n4658, B2 => n10096, C1 => n4722, C2 => 
                           n10092, A => n7844, ZN => n7839);
   U8808 : AOI221_X1 port map( B1 => n4690, B2 => n10112, C1 => n9265, C2 => 
                           n10108, A => n7843, ZN => n7840);
   U8809 : NAND4_X1 port map( A1 => n7821, A2 => n7822, A3 => n7823, A4 => 
                           n7824, ZN => n2358);
   U8810 : AOI221_X1 port map( B1 => n10128, B2 => n7610, C1 => n9330, C2 => 
                           n10124, A => n7825, ZN => n7824);
   U8811 : AOI221_X1 port map( B1 => n4657, B2 => n10096, C1 => n4721, C2 => 
                           n10092, A => n7827, ZN => n7822);
   U8812 : AOI221_X1 port map( B1 => n4689, B2 => n10112, C1 => n9266, C2 => 
                           n10108, A => n7826, ZN => n7823);
   U8813 : NAND4_X1 port map( A1 => n7804, A2 => n7805, A3 => n7806, A4 => 
                           n7807, ZN => n2359);
   U8814 : AOI221_X1 port map( B1 => n10128, B2 => n7609, C1 => n9331, C2 => 
                           n10124, A => n7808, ZN => n7807);
   U8815 : AOI221_X1 port map( B1 => n4656, B2 => n10096, C1 => n4720, C2 => 
                           n10092, A => n7810, ZN => n7805);
   U8816 : AOI221_X1 port map( B1 => n4688, B2 => n10112, C1 => n9267, C2 => 
                           n10108, A => n7809, ZN => n7806);
   U8817 : NAND4_X1 port map( A1 => n7787, A2 => n7788, A3 => n7789, A4 => 
                           n7790, ZN => n2360);
   U8818 : AOI221_X1 port map( B1 => n10129, B2 => n7520, C1 => n9332, C2 => 
                           n10125, A => n7791, ZN => n7790);
   U8819 : AOI221_X1 port map( B1 => n4655, B2 => n10097, C1 => n4719, C2 => 
                           n10093, A => n7793, ZN => n7788);
   U8820 : AOI221_X1 port map( B1 => n4687, B2 => n10113, C1 => n9268, C2 => 
                           n10109, A => n7792, ZN => n7789);
   U8821 : NAND4_X1 port map( A1 => n7770, A2 => n7771, A3 => n7772, A4 => 
                           n7773, ZN => n2361);
   U8822 : AOI221_X1 port map( B1 => n10129, B2 => n7519, C1 => n9333, C2 => 
                           n10125, A => n7774, ZN => n7773);
   U8823 : AOI221_X1 port map( B1 => n4654, B2 => n10097, C1 => n4718, C2 => 
                           n10093, A => n7776, ZN => n7771);
   U8824 : AOI221_X1 port map( B1 => n4686, B2 => n10113, C1 => n9269, C2 => 
                           n10109, A => n7775, ZN => n7772);
   U8825 : NAND4_X1 port map( A1 => n7753, A2 => n7754, A3 => n7755, A4 => 
                           n7756, ZN => n2362);
   U8826 : AOI221_X1 port map( B1 => n10129, B2 => n7518, C1 => n9334, C2 => 
                           n10125, A => n7757, ZN => n7756);
   U8827 : AOI221_X1 port map( B1 => n4653, B2 => n10097, C1 => n4717, C2 => 
                           n10093, A => n7759, ZN => n7754);
   U8828 : AOI221_X1 port map( B1 => n4685, B2 => n10113, C1 => n9270, C2 => 
                           n10109, A => n7758, ZN => n7755);
   U8829 : NAND4_X1 port map( A1 => n7736, A2 => n7737, A3 => n7738, A4 => 
                           n7739, ZN => n2363);
   U8830 : AOI221_X1 port map( B1 => n10129, B2 => n7517, C1 => n9335, C2 => 
                           n10125, A => n7740, ZN => n7739);
   U8831 : AOI221_X1 port map( B1 => n4652, B2 => n10097, C1 => n4716, C2 => 
                           n10093, A => n7742, ZN => n7737);
   U8832 : AOI221_X1 port map( B1 => n4684, B2 => n10113, C1 => n9271, C2 => 
                           n10109, A => n7741, ZN => n7738);
   U8833 : NAND4_X1 port map( A1 => n7719, A2 => n7720, A3 => n7721, A4 => 
                           n7722, ZN => n2364);
   U8834 : AOI221_X1 port map( B1 => n10129, B2 => n7516, C1 => n9336, C2 => 
                           n10125, A => n7723, ZN => n7722);
   U8835 : AOI221_X1 port map( B1 => n4651, B2 => n10097, C1 => n4715, C2 => 
                           n10093, A => n7725, ZN => n7720);
   U8836 : AOI221_X1 port map( B1 => n4683, B2 => n10113, C1 => n9272, C2 => 
                           n10109, A => n7724, ZN => n7721);
   U8837 : NAND4_X1 port map( A1 => n7702, A2 => n7703, A3 => n7704, A4 => 
                           n7705, ZN => n2365);
   U8838 : AOI221_X1 port map( B1 => n10129, B2 => n7515, C1 => n9337, C2 => 
                           n10125, A => n7706, ZN => n7705);
   U8839 : AOI221_X1 port map( B1 => n4650, B2 => n10097, C1 => n4714, C2 => 
                           n10093, A => n7708, ZN => n7703);
   U8840 : AOI221_X1 port map( B1 => n4682, B2 => n10113, C1 => n9273, C2 => 
                           n10109, A => n7707, ZN => n7704);
   U8841 : NAND4_X1 port map( A1 => n7685, A2 => n7686, A3 => n7687, A4 => 
                           n7688, ZN => n2366);
   U8842 : AOI221_X1 port map( B1 => n10129, B2 => n7514, C1 => n9338, C2 => 
                           n10125, A => n7689, ZN => n7688);
   U8843 : AOI221_X1 port map( B1 => n4649, B2 => n10097, C1 => n4713, C2 => 
                           n10093, A => n7691, ZN => n7686);
   U8844 : AOI221_X1 port map( B1 => n4681, B2 => n10113, C1 => n9274, C2 => 
                           n10109, A => n7690, ZN => n7687);
   U8845 : NAND4_X1 port map( A1 => n7634, A2 => n7635, A3 => n7636, A4 => 
                           n7637, ZN => n2367);
   U8846 : AOI221_X1 port map( B1 => n10129, B2 => n7513, C1 => n9339, C2 => 
                           n10125, A => n7640, ZN => n7637);
   U8847 : AOI221_X1 port map( B1 => n4648, B2 => n10097, C1 => n4712, C2 => 
                           n10093, A => n7650, ZN => n7635);
   U8848 : AOI221_X1 port map( B1 => n4680, B2 => n10113, C1 => n9275, C2 => 
                           n10109, A => n7645, ZN => n7636);
   U8849 : AOI221_X1 port map( B1 => n9667, B2 => n9340, C1 => n9663, C2 => 
                           n9180, A => n8886, ZN => n8885);
   U8850 : OAI222_X1 port map( A1 => n7233, A2 => n9659, B1 => n6977, B2 => 
                           n9655, C1 => n7041, C2 => n9651, ZN => n8886);
   U8851 : AOI221_X1 port map( B1 => n9667, B2 => n9341, C1 => n9663, C2 => 
                           n9181, A => n8859, ZN => n8858);
   U8852 : OAI222_X1 port map( A1 => n7232, A2 => n9659, B1 => n6976, B2 => 
                           n9655, C1 => n7040, C2 => n9651, ZN => n8859);
   U8853 : AOI221_X1 port map( B1 => n9667, B2 => n9342, C1 => n9663, C2 => 
                           n9182, A => n8842, ZN => n8841);
   U8854 : OAI222_X1 port map( A1 => n7231, A2 => n9659, B1 => n6975, B2 => 
                           n9655, C1 => n7039, C2 => n9651, ZN => n8842);
   U8855 : AOI221_X1 port map( B1 => n9667, B2 => n9343, C1 => n9663, C2 => 
                           n9183, A => n8825, ZN => n8824);
   U8856 : OAI222_X1 port map( A1 => n7230, A2 => n9659, B1 => n6974, B2 => 
                           n9655, C1 => n7038, C2 => n9651, ZN => n8825);
   U8857 : AOI221_X1 port map( B1 => n9667, B2 => n9344, C1 => n9663, C2 => 
                           n9184, A => n8808, ZN => n8807);
   U8858 : OAI222_X1 port map( A1 => n7229, A2 => n9659, B1 => n6973, B2 => 
                           n9655, C1 => n7037, C2 => n9651, ZN => n8808);
   U8859 : AOI221_X1 port map( B1 => n9667, B2 => n9345, C1 => n9663, C2 => 
                           n9185, A => n8791, ZN => n8790);
   U8860 : OAI222_X1 port map( A1 => n7228, A2 => n9659, B1 => n6972, B2 => 
                           n9655, C1 => n7036, C2 => n9651, ZN => n8791);
   U8861 : AOI221_X1 port map( B1 => n9667, B2 => n9346, C1 => n9663, C2 => 
                           n9186, A => n8774, ZN => n8773);
   U8862 : OAI222_X1 port map( A1 => n7227, A2 => n9659, B1 => n6971, B2 => 
                           n9655, C1 => n7035, C2 => n9651, ZN => n8774);
   U8863 : AOI221_X1 port map( B1 => n9667, B2 => n9347, C1 => n9663, C2 => 
                           n9187, A => n8757, ZN => n8756);
   U8864 : OAI222_X1 port map( A1 => n7226, A2 => n9659, B1 => n6970, B2 => 
                           n9655, C1 => n7034, C2 => n9651, ZN => n8757);
   U8865 : AOI221_X1 port map( B1 => n9667, B2 => n9348, C1 => n9663, C2 => 
                           n9188, A => n8740, ZN => n8739);
   U8866 : OAI222_X1 port map( A1 => n7225, A2 => n9659, B1 => n6969, B2 => 
                           n9655, C1 => n7033, C2 => n9651, ZN => n8740);
   U8867 : AOI221_X1 port map( B1 => n9667, B2 => n9349, C1 => n9663, C2 => 
                           n9189, A => n8723, ZN => n8722);
   U8868 : OAI222_X1 port map( A1 => n7224, A2 => n9659, B1 => n6968, B2 => 
                           n9655, C1 => n7032, C2 => n9651, ZN => n8723);
   U8869 : AOI221_X1 port map( B1 => n9667, B2 => n9350, C1 => n9663, C2 => 
                           n9190, A => n8706, ZN => n8705);
   U8870 : OAI222_X1 port map( A1 => n7223, A2 => n9659, B1 => n6967, B2 => 
                           n9655, C1 => n7031, C2 => n9651, ZN => n8706);
   U8871 : AOI221_X1 port map( B1 => n9667, B2 => n9351, C1 => n9663, C2 => 
                           n9191, A => n8689, ZN => n8688);
   U8872 : OAI222_X1 port map( A1 => n7222, A2 => n9659, B1 => n6966, B2 => 
                           n9655, C1 => n7030, C2 => n9651, ZN => n8689);
   U8873 : AOI221_X1 port map( B1 => n9668, B2 => n9352, C1 => n9664, C2 => 
                           n9192, A => n8672, ZN => n8671);
   U8874 : OAI222_X1 port map( A1 => n7221, A2 => n9660, B1 => n6965, B2 => 
                           n9656, C1 => n7029, C2 => n9652, ZN => n8672);
   U8875 : AOI221_X1 port map( B1 => n9668, B2 => n9353, C1 => n9664, C2 => 
                           n9193, A => n8655, ZN => n8654);
   U8876 : OAI222_X1 port map( A1 => n7220, A2 => n9660, B1 => n6964, B2 => 
                           n9656, C1 => n7028, C2 => n9652, ZN => n8655);
   U8877 : AOI221_X1 port map( B1 => n9668, B2 => n9354, C1 => n9664, C2 => 
                           n9194, A => n8638, ZN => n8637);
   U8878 : OAI222_X1 port map( A1 => n7219, A2 => n9660, B1 => n6963, B2 => 
                           n9656, C1 => n7027, C2 => n9652, ZN => n8638);
   U8879 : AOI221_X1 port map( B1 => n9668, B2 => n9355, C1 => n9664, C2 => 
                           n9195, A => n8621, ZN => n8620);
   U8880 : OAI222_X1 port map( A1 => n7218, A2 => n9660, B1 => n6962, B2 => 
                           n9656, C1 => n7026, C2 => n9652, ZN => n8621);
   U8881 : AOI221_X1 port map( B1 => n9668, B2 => n9356, C1 => n9664, C2 => 
                           n9196, A => n8604, ZN => n8603);
   U8882 : OAI222_X1 port map( A1 => n7217, A2 => n9660, B1 => n6961, B2 => 
                           n9656, C1 => n7025, C2 => n9652, ZN => n8604);
   U8883 : AOI221_X1 port map( B1 => n9668, B2 => n9357, C1 => n9664, C2 => 
                           n9197, A => n8587, ZN => n8586);
   U8884 : OAI222_X1 port map( A1 => n7216, A2 => n9660, B1 => n6960, B2 => 
                           n9656, C1 => n7024, C2 => n9652, ZN => n8587);
   U8885 : AOI221_X1 port map( B1 => n9668, B2 => n9358, C1 => n9664, C2 => 
                           n9198, A => n8570, ZN => n8569);
   U8886 : OAI222_X1 port map( A1 => n7215, A2 => n9660, B1 => n6959, B2 => 
                           n9656, C1 => n7023, C2 => n9652, ZN => n8570);
   U8887 : AOI221_X1 port map( B1 => n9668, B2 => n9359, C1 => n9664, C2 => 
                           n9199, A => n8553, ZN => n8552);
   U8888 : OAI222_X1 port map( A1 => n7214, A2 => n9660, B1 => n6958, B2 => 
                           n9656, C1 => n7022, C2 => n9652, ZN => n8553);
   U8889 : AOI221_X1 port map( B1 => n9668, B2 => n9360, C1 => n9664, C2 => 
                           n9200, A => n8536, ZN => n8535);
   U8890 : OAI222_X1 port map( A1 => n7213, A2 => n9660, B1 => n6957, B2 => 
                           n9656, C1 => n7021, C2 => n9652, ZN => n8536);
   U8891 : AOI221_X1 port map( B1 => n9668, B2 => n9361, C1 => n9664, C2 => 
                           n9201, A => n8519, ZN => n8518);
   U8892 : OAI222_X1 port map( A1 => n7212, A2 => n9660, B1 => n6956, B2 => 
                           n9656, C1 => n7020, C2 => n9652, ZN => n8519);
   U8893 : AOI221_X1 port map( B1 => n9668, B2 => n9362, C1 => n9664, C2 => 
                           n9202, A => n8502, ZN => n8501);
   U8894 : OAI222_X1 port map( A1 => n7211, A2 => n9660, B1 => n6955, B2 => 
                           n9656, C1 => n7019, C2 => n9652, ZN => n8502);
   U8895 : AOI221_X1 port map( B1 => n9668, B2 => n9363, C1 => n9664, C2 => 
                           n9203, A => n8485, ZN => n8484);
   U8896 : OAI222_X1 port map( A1 => n7210, A2 => n9660, B1 => n6954, B2 => 
                           n9656, C1 => n7018, C2 => n9652, ZN => n8485);
   U8897 : AOI221_X1 port map( B1 => n9669, B2 => n9364, C1 => n9665, C2 => 
                           n9204, A => n8468, ZN => n8467);
   U8898 : OAI222_X1 port map( A1 => n7209, A2 => n9661, B1 => n6953, B2 => 
                           n9657, C1 => n7017, C2 => n9653, ZN => n8468);
   U8899 : AOI221_X1 port map( B1 => n9669, B2 => n9365, C1 => n9665, C2 => 
                           n9205, A => n8451, ZN => n8450);
   U8900 : OAI222_X1 port map( A1 => n7208, A2 => n9661, B1 => n6952, B2 => 
                           n9657, C1 => n7016, C2 => n9653, ZN => n8451);
   U8901 : AOI221_X1 port map( B1 => n9669, B2 => n9366, C1 => n9665, C2 => 
                           n9206, A => n8434, ZN => n8433);
   U8902 : OAI222_X1 port map( A1 => n7207, A2 => n9661, B1 => n6951, B2 => 
                           n9657, C1 => n7015, C2 => n9653, ZN => n8434);
   U8903 : AOI221_X1 port map( B1 => n9669, B2 => n9367, C1 => n9665, C2 => 
                           n9207, A => n8417, ZN => n8416);
   U8904 : OAI222_X1 port map( A1 => n7206, A2 => n9661, B1 => n6950, B2 => 
                           n9657, C1 => n7014, C2 => n9653, ZN => n8417);
   U8905 : AOI221_X1 port map( B1 => n9669, B2 => n9368, C1 => n9665, C2 => 
                           n9208, A => n8400, ZN => n8399);
   U8906 : OAI222_X1 port map( A1 => n7205, A2 => n9661, B1 => n6949, B2 => 
                           n9657, C1 => n7013, C2 => n9653, ZN => n8400);
   U8907 : AOI221_X1 port map( B1 => n9669, B2 => n9369, C1 => n9665, C2 => 
                           n9209, A => n8383, ZN => n8382);
   U8908 : OAI222_X1 port map( A1 => n7204, A2 => n9661, B1 => n6948, B2 => 
                           n9657, C1 => n7012, C2 => n9653, ZN => n8383);
   U8909 : AOI221_X1 port map( B1 => n9669, B2 => n9370, C1 => n9665, C2 => 
                           n9210, A => n8366, ZN => n8365);
   U8910 : OAI222_X1 port map( A1 => n7203, A2 => n9661, B1 => n6947, B2 => 
                           n9657, C1 => n7011, C2 => n9653, ZN => n8366);
   U8911 : AOI221_X1 port map( B1 => n9669, B2 => n9371, C1 => n9665, C2 => 
                           n9211, A => n8333, ZN => n8330);
   U8912 : OAI222_X1 port map( A1 => n7202, A2 => n9661, B1 => n6946, B2 => 
                           n9657, C1 => n7010, C2 => n9653, ZN => n8333);
   U8913 : AOI221_X1 port map( B1 => n9684, B2 => n8880, C1 => n9678, C2 => 
                           OUT1_0_port, A => n8881, ZN => n8863);
   U8914 : OAI22_X1 port map( A1 => n7456, A2 => n9674, B1 => n7424, B2 => 
                           n9670, ZN => n8881);
   U8915 : NAND4_X1 port map( A1 => n8882, A2 => n8883, A3 => n8884, A4 => 
                           n8885, ZN => n8880);
   U8916 : AOI221_X1 port map( B1 => n9611, B2 => n9148, C1 => n9607, C2 => 
                           n9020, A => n8891, ZN => n8882);
   U8917 : AOI221_X1 port map( B1 => n9686, B2 => n8853, C1 => n9678, C2 => 
                           OUT1_1_port, A => n8854, ZN => n8846);
   U8918 : OAI22_X1 port map( A1 => n7455, A2 => n9674, B1 => n7423, B2 => 
                           n9670, ZN => n8854);
   U8919 : NAND4_X1 port map( A1 => n8855, A2 => n8856, A3 => n8857, A4 => 
                           n8858, ZN => n8853);
   U8920 : AOI221_X1 port map( B1 => n9611, B2 => n9149, C1 => n9607, C2 => 
                           n9021, A => n8862, ZN => n8855);
   U8921 : AOI221_X1 port map( B1 => n9686, B2 => n8836, C1 => n9678, C2 => 
                           OUT1_2_port, A => n8837, ZN => n8829);
   U8922 : OAI22_X1 port map( A1 => n7454, A2 => n9674, B1 => n7422, B2 => 
                           n9670, ZN => n8837);
   U8923 : NAND4_X1 port map( A1 => n8838, A2 => n8839, A3 => n8840, A4 => 
                           n8841, ZN => n8836);
   U8924 : AOI221_X1 port map( B1 => n9611, B2 => n9150, C1 => n9607, C2 => 
                           n9022, A => n8845, ZN => n8838);
   U8925 : AOI221_X1 port map( B1 => n9685, B2 => n8819, C1 => n9678, C2 => 
                           OUT1_3_port, A => n8820, ZN => n8812);
   U8926 : OAI22_X1 port map( A1 => n7453, A2 => n9674, B1 => n7421, B2 => 
                           n9670, ZN => n8820);
   U8927 : NAND4_X1 port map( A1 => n8821, A2 => n8822, A3 => n8823, A4 => 
                           n8824, ZN => n8819);
   U8928 : AOI221_X1 port map( B1 => n9611, B2 => n9151, C1 => n9607, C2 => 
                           n9023, A => n8828, ZN => n8821);
   U8929 : AOI221_X1 port map( B1 => n9686, B2 => n8802, C1 => n9678, C2 => 
                           OUT1_4_port, A => n8803, ZN => n8795);
   U8930 : OAI22_X1 port map( A1 => n7452, A2 => n9674, B1 => n7420, B2 => 
                           n9670, ZN => n8803);
   U8931 : NAND4_X1 port map( A1 => n8804, A2 => n8805, A3 => n8806, A4 => 
                           n8807, ZN => n8802);
   U8932 : AOI221_X1 port map( B1 => n9611, B2 => n9152, C1 => n9607, C2 => 
                           n9024, A => n8811, ZN => n8804);
   U8933 : AOI221_X1 port map( B1 => n9686, B2 => n8785, C1 => n9678, C2 => 
                           OUT1_5_port, A => n8786, ZN => n8778);
   U8934 : OAI22_X1 port map( A1 => n7451, A2 => n9674, B1 => n7419, B2 => 
                           n9670, ZN => n8786);
   U8935 : NAND4_X1 port map( A1 => n8787, A2 => n8788, A3 => n8789, A4 => 
                           n8790, ZN => n8785);
   U8936 : AOI221_X1 port map( B1 => n9611, B2 => n9153, C1 => n9607, C2 => 
                           n9025, A => n8794, ZN => n8787);
   U8937 : AOI221_X1 port map( B1 => n9686, B2 => n8768, C1 => n9678, C2 => 
                           OUT1_6_port, A => n8769, ZN => n8761);
   U8938 : OAI22_X1 port map( A1 => n7450, A2 => n9674, B1 => n7418, B2 => 
                           n9670, ZN => n8769);
   U8939 : NAND4_X1 port map( A1 => n8770, A2 => n8771, A3 => n8772, A4 => 
                           n8773, ZN => n8768);
   U8940 : AOI221_X1 port map( B1 => n9611, B2 => n9154, C1 => n9607, C2 => 
                           n9026, A => n8777, ZN => n8770);
   U8941 : AOI221_X1 port map( B1 => n9686, B2 => n8751, C1 => n9678, C2 => 
                           OUT1_7_port, A => n8752, ZN => n8744);
   U8942 : OAI22_X1 port map( A1 => n7449, A2 => n9674, B1 => n7417, B2 => 
                           n9670, ZN => n8752);
   U8943 : NAND4_X1 port map( A1 => n8753, A2 => n8754, A3 => n8755, A4 => 
                           n8756, ZN => n8751);
   U8944 : AOI221_X1 port map( B1 => n9611, B2 => n9155, C1 => n9607, C2 => 
                           n9027, A => n8760, ZN => n8753);
   U8945 : AOI221_X1 port map( B1 => n9686, B2 => n8734, C1 => n9678, C2 => 
                           OUT1_8_port, A => n8735, ZN => n8727);
   U8946 : OAI22_X1 port map( A1 => n7448, A2 => n9674, B1 => n7416, B2 => 
                           n9670, ZN => n8735);
   U8947 : NAND4_X1 port map( A1 => n8736, A2 => n8737, A3 => n8738, A4 => 
                           n8739, ZN => n8734);
   U8948 : AOI221_X1 port map( B1 => n9611, B2 => n9156, C1 => n9607, C2 => 
                           n9028, A => n8743, ZN => n8736);
   U8949 : AOI221_X1 port map( B1 => n9686, B2 => n8717, C1 => n9678, C2 => 
                           OUT1_9_port, A => n8718, ZN => n8710);
   U8950 : OAI22_X1 port map( A1 => n7447, A2 => n9674, B1 => n7415, B2 => 
                           n9670, ZN => n8718);
   U8951 : NAND4_X1 port map( A1 => n8719, A2 => n8720, A3 => n8721, A4 => 
                           n8722, ZN => n8717);
   U8952 : AOI221_X1 port map( B1 => n9611, B2 => n9157, C1 => n9607, C2 => 
                           n9029, A => n8726, ZN => n8719);
   U8953 : AOI221_X1 port map( B1 => n9686, B2 => n8700, C1 => n9678, C2 => 
                           OUT1_10_port, A => n8701, ZN => n8693);
   U8954 : OAI22_X1 port map( A1 => n7446, A2 => n9674, B1 => n7414, B2 => 
                           n9670, ZN => n8701);
   U8955 : NAND4_X1 port map( A1 => n8702, A2 => n8703, A3 => n8704, A4 => 
                           n8705, ZN => n8700);
   U8956 : AOI221_X1 port map( B1 => n9611, B2 => n9158, C1 => n9607, C2 => 
                           n9030, A => n8709, ZN => n8702);
   U8957 : AOI221_X1 port map( B1 => n9685, B2 => n8683, C1 => n9678, C2 => 
                           OUT1_11_port, A => n8684, ZN => n8676);
   U8958 : OAI22_X1 port map( A1 => n7445, A2 => n9674, B1 => n7413, B2 => 
                           n9670, ZN => n8684);
   U8959 : NAND4_X1 port map( A1 => n8685, A2 => n8686, A3 => n8687, A4 => 
                           n8688, ZN => n8683);
   U8960 : AOI221_X1 port map( B1 => n9611, B2 => n9159, C1 => n9607, C2 => 
                           n9031, A => n8692, ZN => n8685);
   U8961 : AOI221_X1 port map( B1 => n9685, B2 => n8666, C1 => n9679, C2 => 
                           OUT1_12_port, A => n8667, ZN => n8659);
   U8962 : OAI22_X1 port map( A1 => n7444, A2 => n9675, B1 => n7412, B2 => 
                           n9671, ZN => n8667);
   U8963 : NAND4_X1 port map( A1 => n8668, A2 => n8669, A3 => n8670, A4 => 
                           n8671, ZN => n8666);
   U8964 : AOI221_X1 port map( B1 => n9612, B2 => n9160, C1 => n9608, C2 => 
                           n9032, A => n8675, ZN => n8668);
   U8965 : AOI221_X1 port map( B1 => n9685, B2 => n8649, C1 => n9679, C2 => 
                           OUT1_13_port, A => n8650, ZN => n8642);
   U8966 : OAI22_X1 port map( A1 => n7443, A2 => n9675, B1 => n7411, B2 => 
                           n9671, ZN => n8650);
   U8967 : NAND4_X1 port map( A1 => n8651, A2 => n8652, A3 => n8653, A4 => 
                           n8654, ZN => n8649);
   U8968 : AOI221_X1 port map( B1 => n9612, B2 => n9161, C1 => n9608, C2 => 
                           n9033, A => n8658, ZN => n8651);
   U8969 : AOI221_X1 port map( B1 => n9685, B2 => n8632, C1 => n9679, C2 => 
                           OUT1_14_port, A => n8633, ZN => n8625);
   U8970 : OAI22_X1 port map( A1 => n7442, A2 => n9675, B1 => n7410, B2 => 
                           n9671, ZN => n8633);
   U8971 : NAND4_X1 port map( A1 => n8634, A2 => n8635, A3 => n8636, A4 => 
                           n8637, ZN => n8632);
   U8972 : AOI221_X1 port map( B1 => n9612, B2 => n9162, C1 => n9608, C2 => 
                           n9034, A => n8641, ZN => n8634);
   U8973 : AOI221_X1 port map( B1 => n9685, B2 => n8615, C1 => n9679, C2 => 
                           OUT1_15_port, A => n8616, ZN => n8608);
   U8974 : OAI22_X1 port map( A1 => n7441, A2 => n9675, B1 => n7409, B2 => 
                           n9671, ZN => n8616);
   U8975 : NAND4_X1 port map( A1 => n8617, A2 => n8618, A3 => n8619, A4 => 
                           n8620, ZN => n8615);
   U8976 : AOI221_X1 port map( B1 => n9612, B2 => n9163, C1 => n9608, C2 => 
                           n9035, A => n8624, ZN => n8617);
   U8977 : AOI221_X1 port map( B1 => n9685, B2 => n8598, C1 => n9679, C2 => 
                           OUT1_16_port, A => n8599, ZN => n8591);
   U8978 : OAI22_X1 port map( A1 => n7440, A2 => n9675, B1 => n7408, B2 => 
                           n9671, ZN => n8599);
   U8979 : NAND4_X1 port map( A1 => n8600, A2 => n8601, A3 => n8602, A4 => 
                           n8603, ZN => n8598);
   U8980 : AOI221_X1 port map( B1 => n9612, B2 => n9164, C1 => n9608, C2 => 
                           n9036, A => n8607, ZN => n8600);
   U8981 : AOI221_X1 port map( B1 => n9685, B2 => n8581, C1 => n9679, C2 => 
                           OUT1_17_port, A => n8582, ZN => n8574);
   U8982 : OAI22_X1 port map( A1 => n7439, A2 => n9675, B1 => n7407, B2 => 
                           n9671, ZN => n8582);
   U8983 : NAND4_X1 port map( A1 => n8583, A2 => n8584, A3 => n8585, A4 => 
                           n8586, ZN => n8581);
   U8984 : AOI221_X1 port map( B1 => n9612, B2 => n9165, C1 => n9608, C2 => 
                           n9037, A => n8590, ZN => n8583);
   U8985 : AOI221_X1 port map( B1 => n9685, B2 => n8564, C1 => n9679, C2 => 
                           OUT1_18_port, A => n8565, ZN => n8557);
   U8986 : OAI22_X1 port map( A1 => n7438, A2 => n9675, B1 => n7406, B2 => 
                           n9671, ZN => n8565);
   U8987 : NAND4_X1 port map( A1 => n8566, A2 => n8567, A3 => n8568, A4 => 
                           n8569, ZN => n8564);
   U8988 : AOI221_X1 port map( B1 => n9612, B2 => n9166, C1 => n9608, C2 => 
                           n9038, A => n8573, ZN => n8566);
   U8989 : AOI221_X1 port map( B1 => n9685, B2 => n8547, C1 => n9679, C2 => 
                           OUT1_19_port, A => n8548, ZN => n8540);
   U8990 : OAI22_X1 port map( A1 => n7437, A2 => n9675, B1 => n7405, B2 => 
                           n9671, ZN => n8548);
   U8991 : NAND4_X1 port map( A1 => n8549, A2 => n8550, A3 => n8551, A4 => 
                           n8552, ZN => n8547);
   U8992 : AOI221_X1 port map( B1 => n9612, B2 => n9167, C1 => n9608, C2 => 
                           n9039, A => n8556, ZN => n8549);
   U8993 : AOI221_X1 port map( B1 => n9685, B2 => n8530, C1 => n9679, C2 => 
                           OUT1_20_port, A => n8531, ZN => n8523);
   U8994 : OAI22_X1 port map( A1 => n7436, A2 => n9675, B1 => n7404, B2 => 
                           n9671, ZN => n8531);
   U8995 : NAND4_X1 port map( A1 => n8532, A2 => n8533, A3 => n8534, A4 => 
                           n8535, ZN => n8530);
   U8996 : AOI221_X1 port map( B1 => n9612, B2 => n9168, C1 => n9608, C2 => 
                           n9040, A => n8539, ZN => n8532);
   U8997 : AOI221_X1 port map( B1 => n9685, B2 => n8513, C1 => n9679, C2 => 
                           OUT1_21_port, A => n8514, ZN => n8506);
   U8998 : OAI22_X1 port map( A1 => n7435, A2 => n9675, B1 => n7403, B2 => 
                           n9671, ZN => n8514);
   U8999 : NAND4_X1 port map( A1 => n8515, A2 => n8516, A3 => n8517, A4 => 
                           n8518, ZN => n8513);
   U9000 : AOI221_X1 port map( B1 => n9612, B2 => n9169, C1 => n9608, C2 => 
                           n9041, A => n8522, ZN => n8515);
   U9001 : AOI221_X1 port map( B1 => n9684, B2 => n8496, C1 => n9679, C2 => 
                           OUT1_22_port, A => n8497, ZN => n8489);
   U9002 : OAI22_X1 port map( A1 => n7434, A2 => n9675, B1 => n7402, B2 => 
                           n9671, ZN => n8497);
   U9003 : NAND4_X1 port map( A1 => n8498, A2 => n8499, A3 => n8500, A4 => 
                           n8501, ZN => n8496);
   U9004 : AOI221_X1 port map( B1 => n9612, B2 => n9170, C1 => n9608, C2 => 
                           n9042, A => n8505, ZN => n8498);
   U9005 : AOI221_X1 port map( B1 => n9684, B2 => n8479, C1 => n9679, C2 => 
                           OUT1_23_port, A => n8480, ZN => n8472);
   U9006 : OAI22_X1 port map( A1 => n7433, A2 => n9675, B1 => n7401, B2 => 
                           n9671, ZN => n8480);
   U9007 : NAND4_X1 port map( A1 => n8481, A2 => n8482, A3 => n8483, A4 => 
                           n8484, ZN => n8479);
   U9008 : AOI221_X1 port map( B1 => n9612, B2 => n9171, C1 => n9608, C2 => 
                           n9043, A => n8488, ZN => n8481);
   U9009 : AOI221_X1 port map( B1 => n9684, B2 => n8462, C1 => n9680, C2 => 
                           OUT1_24_port, A => n8463, ZN => n8455);
   U9010 : OAI22_X1 port map( A1 => n7432, A2 => n9676, B1 => n7400, B2 => 
                           n9672, ZN => n8463);
   U9011 : NAND4_X1 port map( A1 => n8464, A2 => n8465, A3 => n8466, A4 => 
                           n8467, ZN => n8462);
   U9012 : AOI221_X1 port map( B1 => n9613, B2 => n9172, C1 => n9609, C2 => 
                           n9044, A => n8471, ZN => n8464);
   U9013 : AOI221_X1 port map( B1 => n9684, B2 => n8445, C1 => n9680, C2 => 
                           OUT1_25_port, A => n8446, ZN => n8438);
   U9014 : OAI22_X1 port map( A1 => n7431, A2 => n9676, B1 => n7399, B2 => 
                           n9672, ZN => n8446);
   U9015 : NAND4_X1 port map( A1 => n8447, A2 => n8448, A3 => n8449, A4 => 
                           n8450, ZN => n8445);
   U9016 : AOI221_X1 port map( B1 => n9613, B2 => n9173, C1 => n9609, C2 => 
                           n9045, A => n8454, ZN => n8447);
   U9017 : AOI221_X1 port map( B1 => n9684, B2 => n8428, C1 => n9680, C2 => 
                           OUT1_26_port, A => n8429, ZN => n8421);
   U9018 : OAI22_X1 port map( A1 => n7430, A2 => n9676, B1 => n7398, B2 => 
                           n9672, ZN => n8429);
   U9019 : NAND4_X1 port map( A1 => n8430, A2 => n8431, A3 => n8432, A4 => 
                           n8433, ZN => n8428);
   U9020 : AOI221_X1 port map( B1 => n9613, B2 => n9174, C1 => n9609, C2 => 
                           n9046, A => n8437, ZN => n8430);
   U9021 : AOI221_X1 port map( B1 => n9684, B2 => n8411, C1 => n9680, C2 => 
                           OUT1_27_port, A => n8412, ZN => n8404);
   U9022 : OAI22_X1 port map( A1 => n7429, A2 => n9676, B1 => n7397, B2 => 
                           n9672, ZN => n8412);
   U9023 : NAND4_X1 port map( A1 => n8413, A2 => n8414, A3 => n8415, A4 => 
                           n8416, ZN => n8411);
   U9024 : AOI221_X1 port map( B1 => n9613, B2 => n9175, C1 => n9609, C2 => 
                           n9047, A => n8420, ZN => n8413);
   U9025 : AOI221_X1 port map( B1 => n9684, B2 => n8394, C1 => n9680, C2 => 
                           OUT1_28_port, A => n8395, ZN => n8387);
   U9026 : OAI22_X1 port map( A1 => n7428, A2 => n9676, B1 => n7396, B2 => 
                           n9672, ZN => n8395);
   U9027 : NAND4_X1 port map( A1 => n8396, A2 => n8397, A3 => n8398, A4 => 
                           n8399, ZN => n8394);
   U9028 : AOI221_X1 port map( B1 => n9613, B2 => n9176, C1 => n9609, C2 => 
                           n9048, A => n8403, ZN => n8396);
   U9029 : AOI221_X1 port map( B1 => n9684, B2 => n8377, C1 => n9680, C2 => 
                           OUT1_29_port, A => n8378, ZN => n8370);
   U9030 : OAI22_X1 port map( A1 => n7427, A2 => n9676, B1 => n7395, B2 => 
                           n9672, ZN => n8378);
   U9031 : NAND4_X1 port map( A1 => n8379, A2 => n8380, A3 => n8381, A4 => 
                           n8382, ZN => n8377);
   U9032 : AOI221_X1 port map( B1 => n9613, B2 => n9177, C1 => n9609, C2 => 
                           n9049, A => n8386, ZN => n8379);
   U9033 : AOI221_X1 port map( B1 => n9684, B2 => n8360, C1 => n9680, C2 => 
                           OUT1_30_port, A => n8361, ZN => n8353);
   U9034 : OAI22_X1 port map( A1 => n7426, A2 => n9676, B1 => n7394, B2 => 
                           n9672, ZN => n8361);
   U9035 : NAND4_X1 port map( A1 => n8362, A2 => n8363, A3 => n8364, A4 => 
                           n8365, ZN => n8360);
   U9036 : AOI221_X1 port map( B1 => n9613, B2 => n9178, C1 => n9609, C2 => 
                           n9050, A => n8369, ZN => n8362);
   U9037 : AOI221_X1 port map( B1 => n9684, B2 => n8322, C1 => n9680, C2 => 
                           OUT1_31_port, A => n8324, ZN => n8302);
   U9038 : OAI22_X1 port map( A1 => n7425, A2 => n9676, B1 => n7393, B2 => 
                           n9672, ZN => n8324);
   U9039 : NAND4_X1 port map( A1 => n8327, A2 => n8328, A3 => n8329, A4 => 
                           n8330, ZN => n8322);
   U9040 : AOI221_X1 port map( B1 => n9613, B2 => n9179, C1 => n9609, C2 => 
                           n9051, A => n8350, ZN => n8327);
   U9041 : NAND4_X1 port map( A1 => n8863, A2 => n8864, A3 => n8865, A4 => 
                           n8866, ZN => n1280);
   U9042 : AOI221_X1 port map( B1 => n9733, B2 => n7632, C1 => n9729, C2 => 
                           n9308, A => n8867, ZN => n8866);
   U9043 : AOI221_X1 port map( B1 => n9701, B2 => n4679, C1 => n9697, C2 => 
                           n4743, A => n8879, ZN => n8864);
   U9044 : AOI221_X1 port map( B1 => n9717, B2 => n4711, C1 => n9713, C2 => 
                           n9244, A => n8873, ZN => n8865);
   U9045 : NAND4_X1 port map( A1 => n8846, A2 => n8847, A3 => n8848, A4 => 
                           n8849, ZN => n1281);
   U9046 : AOI221_X1 port map( B1 => n9733, B2 => n7631, C1 => n9729, C2 => 
                           n9309, A => n8850, ZN => n8849);
   U9047 : AOI221_X1 port map( B1 => n9701, B2 => n4678, C1 => n9697, C2 => 
                           n4742, A => n8852, ZN => n8847);
   U9048 : AOI221_X1 port map( B1 => n9717, B2 => n4710, C1 => n9713, C2 => 
                           n9245, A => n8851, ZN => n8848);
   U9049 : NAND4_X1 port map( A1 => n8829, A2 => n8830, A3 => n8831, A4 => 
                           n8832, ZN => n1282);
   U9050 : AOI221_X1 port map( B1 => n9733, B2 => n7630, C1 => n9729, C2 => 
                           n9310, A => n8833, ZN => n8832);
   U9051 : AOI221_X1 port map( B1 => n9701, B2 => n4677, C1 => n9697, C2 => 
                           n4741, A => n8835, ZN => n8830);
   U9052 : AOI221_X1 port map( B1 => n9717, B2 => n4709, C1 => n9713, C2 => 
                           n9246, A => n8834, ZN => n8831);
   U9053 : NAND4_X1 port map( A1 => n8812, A2 => n8813, A3 => n8814, A4 => 
                           n8815, ZN => n1283);
   U9054 : AOI221_X1 port map( B1 => n9733, B2 => n7629, C1 => n9729, C2 => 
                           n9311, A => n8816, ZN => n8815);
   U9055 : AOI221_X1 port map( B1 => n9701, B2 => n4676, C1 => n9697, C2 => 
                           n4740, A => n8818, ZN => n8813);
   U9056 : AOI221_X1 port map( B1 => n9717, B2 => n4708, C1 => n9713, C2 => 
                           n9247, A => n8817, ZN => n8814);
   U9057 : NAND4_X1 port map( A1 => n8795, A2 => n8796, A3 => n8797, A4 => 
                           n8798, ZN => n1284);
   U9058 : AOI221_X1 port map( B1 => n9733, B2 => n7628, C1 => n9729, C2 => 
                           n9312, A => n8799, ZN => n8798);
   U9059 : AOI221_X1 port map( B1 => n9701, B2 => n4675, C1 => n9697, C2 => 
                           n4739, A => n8801, ZN => n8796);
   U9060 : AOI221_X1 port map( B1 => n9717, B2 => n4707, C1 => n9713, C2 => 
                           n9248, A => n8800, ZN => n8797);
   U9061 : NAND4_X1 port map( A1 => n8778, A2 => n8779, A3 => n8780, A4 => 
                           n8781, ZN => n1285);
   U9062 : AOI221_X1 port map( B1 => n9733, B2 => n7627, C1 => n9729, C2 => 
                           n9313, A => n8782, ZN => n8781);
   U9063 : AOI221_X1 port map( B1 => n9701, B2 => n4674, C1 => n9697, C2 => 
                           n4738, A => n8784, ZN => n8779);
   U9064 : AOI221_X1 port map( B1 => n9717, B2 => n4706, C1 => n9713, C2 => 
                           n9249, A => n8783, ZN => n8780);
   U9065 : NAND4_X1 port map( A1 => n8761, A2 => n8762, A3 => n8763, A4 => 
                           n8764, ZN => n1286);
   U9066 : AOI221_X1 port map( B1 => n9733, B2 => n7626, C1 => n9729, C2 => 
                           n9314, A => n8765, ZN => n8764);
   U9067 : AOI221_X1 port map( B1 => n9701, B2 => n4673, C1 => n9697, C2 => 
                           n4737, A => n8767, ZN => n8762);
   U9068 : AOI221_X1 port map( B1 => n9717, B2 => n4705, C1 => n9713, C2 => 
                           n9250, A => n8766, ZN => n8763);
   U9069 : NAND4_X1 port map( A1 => n8744, A2 => n8745, A3 => n8746, A4 => 
                           n8747, ZN => n1287);
   U9070 : AOI221_X1 port map( B1 => n9733, B2 => n7625, C1 => n9729, C2 => 
                           n9315, A => n8748, ZN => n8747);
   U9071 : AOI221_X1 port map( B1 => n9701, B2 => n4672, C1 => n9697, C2 => 
                           n4736, A => n8750, ZN => n8745);
   U9072 : AOI221_X1 port map( B1 => n9717, B2 => n4704, C1 => n9713, C2 => 
                           n9251, A => n8749, ZN => n8746);
   U9073 : NAND4_X1 port map( A1 => n8727, A2 => n8728, A3 => n8729, A4 => 
                           n8730, ZN => n1288);
   U9074 : AOI221_X1 port map( B1 => n9733, B2 => n7624, C1 => n9729, C2 => 
                           n9316, A => n8731, ZN => n8730);
   U9075 : AOI221_X1 port map( B1 => n9701, B2 => n4671, C1 => n9697, C2 => 
                           n4735, A => n8733, ZN => n8728);
   U9076 : AOI221_X1 port map( B1 => n9717, B2 => n4703, C1 => n9713, C2 => 
                           n9252, A => n8732, ZN => n8729);
   U9077 : NAND4_X1 port map( A1 => n8710, A2 => n8711, A3 => n8712, A4 => 
                           n8713, ZN => n1289);
   U9078 : AOI221_X1 port map( B1 => n9733, B2 => n7623, C1 => n9729, C2 => 
                           n9317, A => n8714, ZN => n8713);
   U9079 : AOI221_X1 port map( B1 => n9701, B2 => n4670, C1 => n9697, C2 => 
                           n4734, A => n8716, ZN => n8711);
   U9080 : AOI221_X1 port map( B1 => n9717, B2 => n4702, C1 => n9713, C2 => 
                           n9253, A => n8715, ZN => n8712);
   U9081 : NAND4_X1 port map( A1 => n8693, A2 => n8694, A3 => n8695, A4 => 
                           n8696, ZN => n1290);
   U9082 : AOI221_X1 port map( B1 => n9733, B2 => n7622, C1 => n9729, C2 => 
                           n9318, A => n8697, ZN => n8696);
   U9083 : AOI221_X1 port map( B1 => n9701, B2 => n4669, C1 => n9697, C2 => 
                           n4733, A => n8699, ZN => n8694);
   U9084 : AOI221_X1 port map( B1 => n9717, B2 => n4701, C1 => n9713, C2 => 
                           n9254, A => n8698, ZN => n8695);
   U9085 : NAND4_X1 port map( A1 => n8676, A2 => n8677, A3 => n8678, A4 => 
                           n8679, ZN => n1291);
   U9086 : AOI221_X1 port map( B1 => n9733, B2 => n7621, C1 => n9729, C2 => 
                           n9319, A => n8680, ZN => n8679);
   U9087 : AOI221_X1 port map( B1 => n9701, B2 => n4668, C1 => n9697, C2 => 
                           n4732, A => n8682, ZN => n8677);
   U9088 : AOI221_X1 port map( B1 => n9717, B2 => n4700, C1 => n9713, C2 => 
                           n9255, A => n8681, ZN => n8678);
   U9089 : NAND4_X1 port map( A1 => n8659, A2 => n8660, A3 => n8661, A4 => 
                           n8662, ZN => n1292);
   U9090 : AOI221_X1 port map( B1 => n9734, B2 => n7620, C1 => n9730, C2 => 
                           n9320, A => n8663, ZN => n8662);
   U9091 : AOI221_X1 port map( B1 => n9702, B2 => n4667, C1 => n9698, C2 => 
                           n4731, A => n8665, ZN => n8660);
   U9092 : AOI221_X1 port map( B1 => n9718, B2 => n4699, C1 => n9714, C2 => 
                           n9256, A => n8664, ZN => n8661);
   U9093 : NAND4_X1 port map( A1 => n8642, A2 => n8643, A3 => n8644, A4 => 
                           n8645, ZN => n1293);
   U9094 : AOI221_X1 port map( B1 => n9734, B2 => n7619, C1 => n9730, C2 => 
                           n9321, A => n8646, ZN => n8645);
   U9095 : AOI221_X1 port map( B1 => n9702, B2 => n4666, C1 => n9698, C2 => 
                           n4730, A => n8648, ZN => n8643);
   U9096 : AOI221_X1 port map( B1 => n9718, B2 => n4698, C1 => n9714, C2 => 
                           n9257, A => n8647, ZN => n8644);
   U9097 : NAND4_X1 port map( A1 => n8625, A2 => n8626, A3 => n8627, A4 => 
                           n8628, ZN => n1294);
   U9098 : AOI221_X1 port map( B1 => n9734, B2 => n7618, C1 => n9730, C2 => 
                           n9322, A => n8629, ZN => n8628);
   U9099 : AOI221_X1 port map( B1 => n9702, B2 => n4665, C1 => n9698, C2 => 
                           n4729, A => n8631, ZN => n8626);
   U9100 : AOI221_X1 port map( B1 => n9718, B2 => n4697, C1 => n9714, C2 => 
                           n9258, A => n8630, ZN => n8627);
   U9101 : NAND4_X1 port map( A1 => n8608, A2 => n8609, A3 => n8610, A4 => 
                           n8611, ZN => n1295);
   U9102 : AOI221_X1 port map( B1 => n9734, B2 => n7617, C1 => n9730, C2 => 
                           n9323, A => n8612, ZN => n8611);
   U9103 : AOI221_X1 port map( B1 => n9702, B2 => n4664, C1 => n9698, C2 => 
                           n4728, A => n8614, ZN => n8609);
   U9104 : AOI221_X1 port map( B1 => n9718, B2 => n4696, C1 => n9714, C2 => 
                           n9259, A => n8613, ZN => n8610);
   U9105 : NAND4_X1 port map( A1 => n8591, A2 => n8592, A3 => n8593, A4 => 
                           n8594, ZN => n1296);
   U9106 : AOI221_X1 port map( B1 => n9734, B2 => n7616, C1 => n9730, C2 => 
                           n9324, A => n8595, ZN => n8594);
   U9107 : AOI221_X1 port map( B1 => n9702, B2 => n4663, C1 => n9698, C2 => 
                           n4727, A => n8597, ZN => n8592);
   U9108 : AOI221_X1 port map( B1 => n9718, B2 => n4695, C1 => n9714, C2 => 
                           n9260, A => n8596, ZN => n8593);
   U9109 : NAND4_X1 port map( A1 => n8574, A2 => n8575, A3 => n8576, A4 => 
                           n8577, ZN => n1297);
   U9110 : AOI221_X1 port map( B1 => n9734, B2 => n7615, C1 => n9730, C2 => 
                           n9325, A => n8578, ZN => n8577);
   U9111 : AOI221_X1 port map( B1 => n9702, B2 => n4662, C1 => n9698, C2 => 
                           n4726, A => n8580, ZN => n8575);
   U9112 : AOI221_X1 port map( B1 => n9718, B2 => n4694, C1 => n9714, C2 => 
                           n9261, A => n8579, ZN => n8576);
   U9113 : NAND4_X1 port map( A1 => n8557, A2 => n8558, A3 => n8559, A4 => 
                           n8560, ZN => n1298);
   U9114 : AOI221_X1 port map( B1 => n9734, B2 => n7614, C1 => n9730, C2 => 
                           n9326, A => n8561, ZN => n8560);
   U9115 : AOI221_X1 port map( B1 => n9702, B2 => n4661, C1 => n9698, C2 => 
                           n4725, A => n8563, ZN => n8558);
   U9116 : AOI221_X1 port map( B1 => n9718, B2 => n4693, C1 => n9714, C2 => 
                           n9262, A => n8562, ZN => n8559);
   U9117 : NAND4_X1 port map( A1 => n8540, A2 => n8541, A3 => n8542, A4 => 
                           n8543, ZN => n1299);
   U9118 : AOI221_X1 port map( B1 => n9734, B2 => n7613, C1 => n9730, C2 => 
                           n9327, A => n8544, ZN => n8543);
   U9119 : AOI221_X1 port map( B1 => n9702, B2 => n4660, C1 => n9698, C2 => 
                           n4724, A => n8546, ZN => n8541);
   U9120 : AOI221_X1 port map( B1 => n9718, B2 => n4692, C1 => n9714, C2 => 
                           n9263, A => n8545, ZN => n8542);
   U9121 : NAND4_X1 port map( A1 => n8523, A2 => n8524, A3 => n8525, A4 => 
                           n8526, ZN => n1300);
   U9122 : AOI221_X1 port map( B1 => n9734, B2 => n7612, C1 => n9730, C2 => 
                           n9328, A => n8527, ZN => n8526);
   U9123 : AOI221_X1 port map( B1 => n9702, B2 => n4659, C1 => n9698, C2 => 
                           n4723, A => n8529, ZN => n8524);
   U9124 : AOI221_X1 port map( B1 => n9718, B2 => n4691, C1 => n9714, C2 => 
                           n9264, A => n8528, ZN => n8525);
   U9125 : NAND4_X1 port map( A1 => n8506, A2 => n8507, A3 => n8508, A4 => 
                           n8509, ZN => n1301);
   U9126 : AOI221_X1 port map( B1 => n9734, B2 => n7611, C1 => n9730, C2 => 
                           n9329, A => n8510, ZN => n8509);
   U9127 : AOI221_X1 port map( B1 => n9702, B2 => n4658, C1 => n9698, C2 => 
                           n4722, A => n8512, ZN => n8507);
   U9128 : AOI221_X1 port map( B1 => n9718, B2 => n4690, C1 => n9714, C2 => 
                           n9265, A => n8511, ZN => n8508);
   U9129 : NAND4_X1 port map( A1 => n8489, A2 => n8490, A3 => n8491, A4 => 
                           n8492, ZN => n1302);
   U9130 : AOI221_X1 port map( B1 => n9734, B2 => n7610, C1 => n9730, C2 => 
                           n9330, A => n8493, ZN => n8492);
   U9131 : AOI221_X1 port map( B1 => n9702, B2 => n4657, C1 => n9698, C2 => 
                           n4721, A => n8495, ZN => n8490);
   U9132 : AOI221_X1 port map( B1 => n9718, B2 => n4689, C1 => n9714, C2 => 
                           n9266, A => n8494, ZN => n8491);
   U9133 : NAND4_X1 port map( A1 => n8472, A2 => n8473, A3 => n8474, A4 => 
                           n8475, ZN => n1303);
   U9134 : AOI221_X1 port map( B1 => n9734, B2 => n7609, C1 => n9730, C2 => 
                           n9331, A => n8476, ZN => n8475);
   U9135 : AOI221_X1 port map( B1 => n9702, B2 => n4656, C1 => n9698, C2 => 
                           n4720, A => n8478, ZN => n8473);
   U9136 : AOI221_X1 port map( B1 => n9718, B2 => n4688, C1 => n9714, C2 => 
                           n9267, A => n8477, ZN => n8474);
   U9137 : NAND4_X1 port map( A1 => n8455, A2 => n8456, A3 => n8457, A4 => 
                           n8458, ZN => n1304);
   U9138 : AOI221_X1 port map( B1 => n9735, B2 => n7520, C1 => n9731, C2 => 
                           n9332, A => n8459, ZN => n8458);
   U9139 : AOI221_X1 port map( B1 => n9703, B2 => n4655, C1 => n9699, C2 => 
                           n4719, A => n8461, ZN => n8456);
   U9140 : AOI221_X1 port map( B1 => n9719, B2 => n4687, C1 => n9715, C2 => 
                           n9268, A => n8460, ZN => n8457);
   U9141 : NAND4_X1 port map( A1 => n8438, A2 => n8439, A3 => n8440, A4 => 
                           n8441, ZN => n1305);
   U9142 : AOI221_X1 port map( B1 => n9735, B2 => n7519, C1 => n9731, C2 => 
                           n9333, A => n8442, ZN => n8441);
   U9143 : AOI221_X1 port map( B1 => n9703, B2 => n4654, C1 => n9699, C2 => 
                           n4718, A => n8444, ZN => n8439);
   U9144 : AOI221_X1 port map( B1 => n9719, B2 => n4686, C1 => n9715, C2 => 
                           n9269, A => n8443, ZN => n8440);
   U9145 : NAND4_X1 port map( A1 => n8421, A2 => n8422, A3 => n8423, A4 => 
                           n8424, ZN => n1306);
   U9146 : AOI221_X1 port map( B1 => n9735, B2 => n7518, C1 => n9731, C2 => 
                           n9334, A => n8425, ZN => n8424);
   U9147 : AOI221_X1 port map( B1 => n9703, B2 => n4653, C1 => n9699, C2 => 
                           n4717, A => n8427, ZN => n8422);
   U9148 : AOI221_X1 port map( B1 => n9719, B2 => n4685, C1 => n9715, C2 => 
                           n9270, A => n8426, ZN => n8423);
   U9149 : NAND4_X1 port map( A1 => n8404, A2 => n8405, A3 => n8406, A4 => 
                           n8407, ZN => n1307);
   U9150 : AOI221_X1 port map( B1 => n9735, B2 => n7517, C1 => n9731, C2 => 
                           n9335, A => n8408, ZN => n8407);
   U9151 : AOI221_X1 port map( B1 => n9703, B2 => n4652, C1 => n9699, C2 => 
                           n4716, A => n8410, ZN => n8405);
   U9152 : AOI221_X1 port map( B1 => n9719, B2 => n4684, C1 => n9715, C2 => 
                           n9271, A => n8409, ZN => n8406);
   U9153 : NAND4_X1 port map( A1 => n8387, A2 => n8388, A3 => n8389, A4 => 
                           n8390, ZN => n1308);
   U9154 : AOI221_X1 port map( B1 => n9735, B2 => n7516, C1 => n9731, C2 => 
                           n9336, A => n8391, ZN => n8390);
   U9155 : AOI221_X1 port map( B1 => n9703, B2 => n4651, C1 => n9699, C2 => 
                           n4715, A => n8393, ZN => n8388);
   U9156 : AOI221_X1 port map( B1 => n9719, B2 => n4683, C1 => n9715, C2 => 
                           n9272, A => n8392, ZN => n8389);
   U9157 : NAND4_X1 port map( A1 => n8370, A2 => n8371, A3 => n8372, A4 => 
                           n8373, ZN => n1309);
   U9158 : AOI221_X1 port map( B1 => n9735, B2 => n7515, C1 => n9731, C2 => 
                           n9337, A => n8374, ZN => n8373);
   U9159 : AOI221_X1 port map( B1 => n9703, B2 => n4650, C1 => n9699, C2 => 
                           n4714, A => n8376, ZN => n8371);
   U9160 : AOI221_X1 port map( B1 => n9719, B2 => n4682, C1 => n9715, C2 => 
                           n9273, A => n8375, ZN => n8372);
   U9161 : NAND4_X1 port map( A1 => n8353, A2 => n8354, A3 => n8355, A4 => 
                           n8356, ZN => n1310);
   U9162 : AOI221_X1 port map( B1 => n9735, B2 => n7514, C1 => n9731, C2 => 
                           n9338, A => n8357, ZN => n8356);
   U9163 : AOI221_X1 port map( B1 => n9703, B2 => n4649, C1 => n9699, C2 => 
                           n4713, A => n8359, ZN => n8354);
   U9164 : AOI221_X1 port map( B1 => n9719, B2 => n4681, C1 => n9715, C2 => 
                           n9274, A => n8358, ZN => n8355);
   U9165 : NAND4_X1 port map( A1 => n8302, A2 => n8303, A3 => n8304, A4 => 
                           n8305, ZN => n1311);
   U9166 : AOI221_X1 port map( B1 => n9735, B2 => n7513, C1 => n9731, C2 => 
                           n9339, A => n8308, ZN => n8305);
   U9167 : AOI221_X1 port map( B1 => n9703, B2 => n4648, C1 => n9699, C2 => 
                           n4712, A => n8318, ZN => n8303);
   U9168 : AOI221_X1 port map( B1 => n9719, B2 => n4680, C1 => n9715, C2 => 
                           n9275, A => n8313, ZN => n8304);
   U9169 : AOI221_X1 port map( B1 => n9532, B2 => n10025, C1 => n9404, C2 => 
                           n10021, A => n8222, ZN => n8215);
   U9170 : OAI222_X1 port map( A1 => n10017, A2 => n7009, B1 => n10013, B2 => 
                           n7137, C1 => n10009, C2 => n7265, ZN => n8222);
   U9171 : AOI221_X1 port map( B1 => n9533, B2 => n10025, C1 => n9405, C2 => 
                           n10021, A => n8193, ZN => n8188);
   U9172 : OAI222_X1 port map( A1 => n10017, A2 => n7008, B1 => n10013, B2 => 
                           n7136, C1 => n10009, C2 => n7264, ZN => n8193);
   U9173 : AOI221_X1 port map( B1 => n9534, B2 => n10025, C1 => n9406, C2 => 
                           n10021, A => n8176, ZN => n8171);
   U9174 : OAI222_X1 port map( A1 => n10017, A2 => n7007, B1 => n10013, B2 => 
                           n7135, C1 => n10009, C2 => n7263, ZN => n8176);
   U9175 : AOI221_X1 port map( B1 => n9535, B2 => n10025, C1 => n9407, C2 => 
                           n10021, A => n8159, ZN => n8154);
   U9176 : OAI222_X1 port map( A1 => n10017, A2 => n7006, B1 => n10013, B2 => 
                           n7134, C1 => n10009, C2 => n7262, ZN => n8159);
   U9177 : AOI221_X1 port map( B1 => n9536, B2 => n10025, C1 => n9408, C2 => 
                           n10021, A => n8142, ZN => n8137);
   U9178 : OAI222_X1 port map( A1 => n10017, A2 => n7005, B1 => n10013, B2 => 
                           n7133, C1 => n10009, C2 => n7261, ZN => n8142);
   U9179 : AOI221_X1 port map( B1 => n9537, B2 => n10025, C1 => n9409, C2 => 
                           n10021, A => n8125, ZN => n8120);
   U9180 : OAI222_X1 port map( A1 => n10017, A2 => n7004, B1 => n10013, B2 => 
                           n7132, C1 => n10009, C2 => n7260, ZN => n8125);
   U9181 : AOI221_X1 port map( B1 => n9538, B2 => n10025, C1 => n9410, C2 => 
                           n10021, A => n8108, ZN => n8103);
   U9182 : OAI222_X1 port map( A1 => n10017, A2 => n7003, B1 => n10013, B2 => 
                           n7131, C1 => n10009, C2 => n7259, ZN => n8108);
   U9183 : AOI221_X1 port map( B1 => n9539, B2 => n10025, C1 => n9411, C2 => 
                           n10021, A => n8091, ZN => n8086);
   U9184 : OAI222_X1 port map( A1 => n10017, A2 => n7002, B1 => n10013, B2 => 
                           n7130, C1 => n10009, C2 => n7258, ZN => n8091);
   U9185 : AOI221_X1 port map( B1 => n9540, B2 => n10025, C1 => n9412, C2 => 
                           n10021, A => n8074, ZN => n8069);
   U9186 : OAI222_X1 port map( A1 => n10017, A2 => n7001, B1 => n10013, B2 => 
                           n7129, C1 => n10009, C2 => n7257, ZN => n8074);
   U9187 : AOI221_X1 port map( B1 => n9541, B2 => n10025, C1 => n9413, C2 => 
                           n10021, A => n8057, ZN => n8052);
   U9188 : OAI222_X1 port map( A1 => n10017, A2 => n7000, B1 => n10013, B2 => 
                           n7128, C1 => n10009, C2 => n7256, ZN => n8057);
   U9189 : AOI221_X1 port map( B1 => n9542, B2 => n10025, C1 => n9414, C2 => 
                           n10021, A => n8040, ZN => n8035);
   U9190 : OAI222_X1 port map( A1 => n10017, A2 => n6999, B1 => n10013, B2 => 
                           n7127, C1 => n10009, C2 => n7255, ZN => n8040);
   U9191 : AOI221_X1 port map( B1 => n9543, B2 => n10025, C1 => n9415, C2 => 
                           n10021, A => n8023, ZN => n8018);
   U9192 : OAI222_X1 port map( A1 => n10017, A2 => n6998, B1 => n10013, B2 => 
                           n7126, C1 => n10009, C2 => n7254, ZN => n8023);
   U9193 : AOI221_X1 port map( B1 => n9544, B2 => n10026, C1 => n9416, C2 => 
                           n10022, A => n8006, ZN => n8001);
   U9194 : OAI222_X1 port map( A1 => n10018, A2 => n6997, B1 => n10014, B2 => 
                           n7125, C1 => n10010, C2 => n7253, ZN => n8006);
   U9195 : AOI221_X1 port map( B1 => n9545, B2 => n10026, C1 => n9417, C2 => 
                           n10022, A => n7989, ZN => n7984);
   U9196 : OAI222_X1 port map( A1 => n10018, A2 => n6996, B1 => n10014, B2 => 
                           n7124, C1 => n10010, C2 => n7252, ZN => n7989);
   U9197 : AOI221_X1 port map( B1 => n9546, B2 => n10026, C1 => n9418, C2 => 
                           n10022, A => n7972, ZN => n7967);
   U9198 : OAI222_X1 port map( A1 => n10018, A2 => n6995, B1 => n10014, B2 => 
                           n7123, C1 => n10010, C2 => n7251, ZN => n7972);
   U9199 : AOI221_X1 port map( B1 => n9547, B2 => n10026, C1 => n9419, C2 => 
                           n10022, A => n7955, ZN => n7950);
   U9200 : OAI222_X1 port map( A1 => n10018, A2 => n6994, B1 => n10014, B2 => 
                           n7122, C1 => n10010, C2 => n7250, ZN => n7955);
   U9201 : AOI221_X1 port map( B1 => n9548, B2 => n10026, C1 => n9420, C2 => 
                           n10022, A => n7938, ZN => n7933);
   U9202 : OAI222_X1 port map( A1 => n10018, A2 => n6993, B1 => n10014, B2 => 
                           n7121, C1 => n10010, C2 => n7249, ZN => n7938);
   U9203 : AOI221_X1 port map( B1 => n9549, B2 => n10026, C1 => n9421, C2 => 
                           n10022, A => n7921, ZN => n7916);
   U9204 : OAI222_X1 port map( A1 => n10018, A2 => n6992, B1 => n10014, B2 => 
                           n7120, C1 => n10010, C2 => n7248, ZN => n7921);
   U9205 : AOI221_X1 port map( B1 => n9550, B2 => n10026, C1 => n9422, C2 => 
                           n10022, A => n7904, ZN => n7899);
   U9206 : OAI222_X1 port map( A1 => n10018, A2 => n6991, B1 => n10014, B2 => 
                           n7119, C1 => n10010, C2 => n7247, ZN => n7904);
   U9207 : AOI221_X1 port map( B1 => n9551, B2 => n10026, C1 => n9423, C2 => 
                           n10022, A => n7887, ZN => n7882);
   U9208 : OAI222_X1 port map( A1 => n10018, A2 => n6990, B1 => n10014, B2 => 
                           n7118, C1 => n10010, C2 => n7246, ZN => n7887);
   U9209 : AOI221_X1 port map( B1 => n9552, B2 => n10026, C1 => n9424, C2 => 
                           n10022, A => n7870, ZN => n7865);
   U9210 : OAI222_X1 port map( A1 => n10018, A2 => n6989, B1 => n10014, B2 => 
                           n7117, C1 => n10010, C2 => n7245, ZN => n7870);
   U9211 : AOI221_X1 port map( B1 => n9553, B2 => n10026, C1 => n9425, C2 => 
                           n10022, A => n7853, ZN => n7848);
   U9212 : OAI222_X1 port map( A1 => n10018, A2 => n6988, B1 => n10014, B2 => 
                           n7116, C1 => n10010, C2 => n7244, ZN => n7853);
   U9213 : AOI221_X1 port map( B1 => n9554, B2 => n10026, C1 => n9426, C2 => 
                           n10022, A => n7836, ZN => n7831);
   U9214 : OAI222_X1 port map( A1 => n10018, A2 => n6987, B1 => n10014, B2 => 
                           n7115, C1 => n10010, C2 => n7243, ZN => n7836);
   U9215 : AOI221_X1 port map( B1 => n9555, B2 => n10026, C1 => n9427, C2 => 
                           n10022, A => n7819, ZN => n7814);
   U9216 : OAI222_X1 port map( A1 => n10018, A2 => n6986, B1 => n10014, B2 => 
                           n7114, C1 => n10010, C2 => n7242, ZN => n7819);
   U9217 : AOI221_X1 port map( B1 => n9556, B2 => n10027, C1 => n9428, C2 => 
                           n10023, A => n7802, ZN => n7797);
   U9218 : OAI222_X1 port map( A1 => n10019, A2 => n6985, B1 => n10015, B2 => 
                           n7113, C1 => n10011, C2 => n7241, ZN => n7802);
   U9219 : AOI221_X1 port map( B1 => n9557, B2 => n10027, C1 => n9429, C2 => 
                           n10023, A => n7785, ZN => n7780);
   U9220 : OAI222_X1 port map( A1 => n10019, A2 => n6984, B1 => n10015, B2 => 
                           n7112, C1 => n10011, C2 => n7240, ZN => n7785);
   U9221 : AOI221_X1 port map( B1 => n9558, B2 => n10027, C1 => n9430, C2 => 
                           n10023, A => n7768, ZN => n7763);
   U9222 : OAI222_X1 port map( A1 => n10019, A2 => n6983, B1 => n10015, B2 => 
                           n7111, C1 => n10011, C2 => n7239, ZN => n7768);
   U9223 : AOI221_X1 port map( B1 => n9559, B2 => n10027, C1 => n9431, C2 => 
                           n10023, A => n7751, ZN => n7746);
   U9224 : OAI222_X1 port map( A1 => n10019, A2 => n6982, B1 => n10015, B2 => 
                           n7110, C1 => n10011, C2 => n7238, ZN => n7751);
   U9225 : AOI221_X1 port map( B1 => n9560, B2 => n10027, C1 => n9432, C2 => 
                           n10023, A => n7734, ZN => n7729);
   U9226 : OAI222_X1 port map( A1 => n10019, A2 => n6981, B1 => n10015, B2 => 
                           n7109, C1 => n10011, C2 => n7237, ZN => n7734);
   U9227 : AOI221_X1 port map( B1 => n9561, B2 => n10027, C1 => n9433, C2 => 
                           n10023, A => n7717, ZN => n7712);
   U9228 : OAI222_X1 port map( A1 => n10019, A2 => n6980, B1 => n10015, B2 => 
                           n7108, C1 => n10011, C2 => n7236, ZN => n7717);
   U9229 : AOI221_X1 port map( B1 => n9562, B2 => n10027, C1 => n9434, C2 => 
                           n10023, A => n7700, ZN => n7695);
   U9230 : OAI222_X1 port map( A1 => n10019, A2 => n6979, B1 => n10015, B2 => 
                           n7107, C1 => n10011, C2 => n7235, ZN => n7700);
   U9231 : AOI221_X1 port map( B1 => n9563, B2 => n10027, C1 => n9435, C2 => 
                           n10023, A => n7676, ZN => n7660);
   U9232 : OAI222_X1 port map( A1 => n10019, A2 => n6978, B1 => n10015, B2 => 
                           n7106, C1 => n10011, C2 => n7234, ZN => n7676);
   U9233 : AOI221_X1 port map( B1 => n9633, B2 => n9556, C1 => n9629, C2 => 
                           n9428, A => n8470, ZN => n8465);
   U9234 : OAI222_X1 port map( A1 => n6985, A2 => n9625, B1 => n7113, B2 => 
                           n9621, C1 => n7241, C2 => n9617, ZN => n8470);
   U9235 : AOI221_X1 port map( B1 => n9633, B2 => n9557, C1 => n9629, C2 => 
                           n9429, A => n8453, ZN => n8448);
   U9236 : OAI222_X1 port map( A1 => n6984, A2 => n9625, B1 => n7112, B2 => 
                           n9621, C1 => n7240, C2 => n9617, ZN => n8453);
   U9237 : AOI221_X1 port map( B1 => n9633, B2 => n9558, C1 => n9629, C2 => 
                           n9430, A => n8436, ZN => n8431);
   U9238 : OAI222_X1 port map( A1 => n6983, A2 => n9625, B1 => n7111, B2 => 
                           n9621, C1 => n7239, C2 => n9617, ZN => n8436);
   U9239 : AOI221_X1 port map( B1 => n9633, B2 => n9559, C1 => n9629, C2 => 
                           n9431, A => n8419, ZN => n8414);
   U9240 : OAI222_X1 port map( A1 => n6982, A2 => n9625, B1 => n7110, B2 => 
                           n9621, C1 => n7238, C2 => n9617, ZN => n8419);
   U9241 : AOI221_X1 port map( B1 => n9633, B2 => n9560, C1 => n9629, C2 => 
                           n9432, A => n8402, ZN => n8397);
   U9242 : OAI222_X1 port map( A1 => n6981, A2 => n9625, B1 => n7109, B2 => 
                           n9621, C1 => n7237, C2 => n9617, ZN => n8402);
   U9243 : AOI221_X1 port map( B1 => n9633, B2 => n9561, C1 => n9629, C2 => 
                           n9433, A => n8385, ZN => n8380);
   U9244 : OAI222_X1 port map( A1 => n6980, A2 => n9625, B1 => n7108, B2 => 
                           n9621, C1 => n7236, C2 => n9617, ZN => n8385);
   U9245 : AOI221_X1 port map( B1 => n9633, B2 => n9562, C1 => n9629, C2 => 
                           n9434, A => n8368, ZN => n8363);
   U9246 : OAI222_X1 port map( A1 => n6979, A2 => n9625, B1 => n7107, B2 => 
                           n9621, C1 => n7235, C2 => n9617, ZN => n8368);
   U9247 : AOI221_X1 port map( B1 => n9633, B2 => n9563, C1 => n9629, C2 => 
                           n9435, A => n8344, ZN => n8328);
   U9248 : OAI222_X1 port map( A1 => n6978, A2 => n9625, B1 => n7106, B2 => 
                           n9621, C1 => n7234, C2 => n9617, ZN => n8344);
   U9249 : AOI221_X1 port map( B1 => n9631, B2 => n9532, C1 => n9627, C2 => 
                           n9404, A => n8890, ZN => n8883);
   U9250 : OAI222_X1 port map( A1 => n7009, A2 => n9623, B1 => n7137, B2 => 
                           n9619, C1 => n7265, C2 => n9615, ZN => n8890);
   U9251 : AOI221_X1 port map( B1 => n9631, B2 => n9533, C1 => n9627, C2 => 
                           n9405, A => n8861, ZN => n8856);
   U9252 : OAI222_X1 port map( A1 => n7008, A2 => n9623, B1 => n7136, B2 => 
                           n9619, C1 => n7264, C2 => n9615, ZN => n8861);
   U9253 : AOI221_X1 port map( B1 => n9631, B2 => n9534, C1 => n9627, C2 => 
                           n9406, A => n8844, ZN => n8839);
   U9254 : OAI222_X1 port map( A1 => n7007, A2 => n9623, B1 => n7135, B2 => 
                           n9619, C1 => n7263, C2 => n9615, ZN => n8844);
   U9255 : AOI221_X1 port map( B1 => n9631, B2 => n9535, C1 => n9627, C2 => 
                           n9407, A => n8827, ZN => n8822);
   U9256 : OAI222_X1 port map( A1 => n7006, A2 => n9623, B1 => n7134, B2 => 
                           n9619, C1 => n7262, C2 => n9615, ZN => n8827);
   U9257 : AOI221_X1 port map( B1 => n9631, B2 => n9536, C1 => n9627, C2 => 
                           n9408, A => n8810, ZN => n8805);
   U9258 : OAI222_X1 port map( A1 => n7005, A2 => n9623, B1 => n7133, B2 => 
                           n9619, C1 => n7261, C2 => n9615, ZN => n8810);
   U9259 : AOI221_X1 port map( B1 => n9631, B2 => n9537, C1 => n9627, C2 => 
                           n9409, A => n8793, ZN => n8788);
   U9260 : OAI222_X1 port map( A1 => n7004, A2 => n9623, B1 => n7132, B2 => 
                           n9619, C1 => n7260, C2 => n9615, ZN => n8793);
   U9261 : AOI221_X1 port map( B1 => n9631, B2 => n9538, C1 => n9627, C2 => 
                           n9410, A => n8776, ZN => n8771);
   U9262 : OAI222_X1 port map( A1 => n7003, A2 => n9623, B1 => n7131, B2 => 
                           n9619, C1 => n7259, C2 => n9615, ZN => n8776);
   U9263 : AOI221_X1 port map( B1 => n9631, B2 => n9539, C1 => n9627, C2 => 
                           n9411, A => n8759, ZN => n8754);
   U9264 : OAI222_X1 port map( A1 => n7002, A2 => n9623, B1 => n7130, B2 => 
                           n9619, C1 => n7258, C2 => n9615, ZN => n8759);
   U9265 : AOI221_X1 port map( B1 => n9631, B2 => n9540, C1 => n9627, C2 => 
                           n9412, A => n8742, ZN => n8737);
   U9266 : OAI222_X1 port map( A1 => n7001, A2 => n9623, B1 => n7129, B2 => 
                           n9619, C1 => n7257, C2 => n9615, ZN => n8742);
   U9267 : AOI221_X1 port map( B1 => n9631, B2 => n9541, C1 => n9627, C2 => 
                           n9413, A => n8725, ZN => n8720);
   U9268 : OAI222_X1 port map( A1 => n7000, A2 => n9623, B1 => n7128, B2 => 
                           n9619, C1 => n7256, C2 => n9615, ZN => n8725);
   U9269 : AOI221_X1 port map( B1 => n9631, B2 => n9542, C1 => n9627, C2 => 
                           n9414, A => n8708, ZN => n8703);
   U9270 : OAI222_X1 port map( A1 => n6999, A2 => n9623, B1 => n7127, B2 => 
                           n9619, C1 => n7255, C2 => n9615, ZN => n8708);
   U9271 : AOI221_X1 port map( B1 => n9631, B2 => n9543, C1 => n9627, C2 => 
                           n9415, A => n8691, ZN => n8686);
   U9272 : OAI222_X1 port map( A1 => n6998, A2 => n9623, B1 => n7126, B2 => 
                           n9619, C1 => n7254, C2 => n9615, ZN => n8691);
   U9273 : AOI221_X1 port map( B1 => n9632, B2 => n9544, C1 => n9628, C2 => 
                           n9416, A => n8674, ZN => n8669);
   U9274 : OAI222_X1 port map( A1 => n6997, A2 => n9624, B1 => n7125, B2 => 
                           n9620, C1 => n7253, C2 => n9616, ZN => n8674);
   U9275 : AOI221_X1 port map( B1 => n9632, B2 => n9545, C1 => n9628, C2 => 
                           n9417, A => n8657, ZN => n8652);
   U9276 : OAI222_X1 port map( A1 => n6996, A2 => n9624, B1 => n7124, B2 => 
                           n9620, C1 => n7252, C2 => n9616, ZN => n8657);
   U9277 : AOI221_X1 port map( B1 => n9632, B2 => n9546, C1 => n9628, C2 => 
                           n9418, A => n8640, ZN => n8635);
   U9278 : OAI222_X1 port map( A1 => n6995, A2 => n9624, B1 => n7123, B2 => 
                           n9620, C1 => n7251, C2 => n9616, ZN => n8640);
   U9279 : AOI221_X1 port map( B1 => n9632, B2 => n9547, C1 => n9628, C2 => 
                           n9419, A => n8623, ZN => n8618);
   U9280 : OAI222_X1 port map( A1 => n6994, A2 => n9624, B1 => n7122, B2 => 
                           n9620, C1 => n7250, C2 => n9616, ZN => n8623);
   U9281 : AOI221_X1 port map( B1 => n9632, B2 => n9548, C1 => n9628, C2 => 
                           n9420, A => n8606, ZN => n8601);
   U9282 : OAI222_X1 port map( A1 => n6993, A2 => n9624, B1 => n7121, B2 => 
                           n9620, C1 => n7249, C2 => n9616, ZN => n8606);
   U9283 : AOI221_X1 port map( B1 => n9632, B2 => n9549, C1 => n9628, C2 => 
                           n9421, A => n8589, ZN => n8584);
   U9284 : OAI222_X1 port map( A1 => n6992, A2 => n9624, B1 => n7120, B2 => 
                           n9620, C1 => n7248, C2 => n9616, ZN => n8589);
   U9285 : AOI221_X1 port map( B1 => n9632, B2 => n9550, C1 => n9628, C2 => 
                           n9422, A => n8572, ZN => n8567);
   U9286 : OAI222_X1 port map( A1 => n6991, A2 => n9624, B1 => n7119, B2 => 
                           n9620, C1 => n7247, C2 => n9616, ZN => n8572);
   U9287 : AOI221_X1 port map( B1 => n9632, B2 => n9551, C1 => n9628, C2 => 
                           n9423, A => n8555, ZN => n8550);
   U9288 : OAI222_X1 port map( A1 => n6990, A2 => n9624, B1 => n7118, B2 => 
                           n9620, C1 => n7246, C2 => n9616, ZN => n8555);
   U9289 : AOI221_X1 port map( B1 => n9632, B2 => n9552, C1 => n9628, C2 => 
                           n9424, A => n8538, ZN => n8533);
   U9290 : OAI222_X1 port map( A1 => n6989, A2 => n9624, B1 => n7117, B2 => 
                           n9620, C1 => n7245, C2 => n9616, ZN => n8538);
   U9291 : AOI221_X1 port map( B1 => n9632, B2 => n9553, C1 => n9628, C2 => 
                           n9425, A => n8521, ZN => n8516);
   U9292 : OAI222_X1 port map( A1 => n6988, A2 => n9624, B1 => n7116, B2 => 
                           n9620, C1 => n7244, C2 => n9616, ZN => n8521);
   U9293 : AOI221_X1 port map( B1 => n9632, B2 => n9554, C1 => n9628, C2 => 
                           n9426, A => n8504, ZN => n8499);
   U9294 : OAI222_X1 port map( A1 => n6987, A2 => n9624, B1 => n7115, B2 => 
                           n9620, C1 => n7243, C2 => n9616, ZN => n8504);
   U9295 : AOI221_X1 port map( B1 => n9632, B2 => n9555, C1 => n9628, C2 => 
                           n9427, A => n8487, ZN => n8482);
   U9296 : OAI222_X1 port map( A1 => n6986, A2 => n9624, B1 => n7114, B2 => 
                           n9620, C1 => n7242, C2 => n9616, ZN => n8487);
   U9297 : AOI221_X1 port map( B1 => n9084, B2 => n10041, C1 => n9564, C2 => 
                           n10037, A => n8221, ZN => n8216);
   U9298 : OAI22_X1 port map( A1 => n10033, A2 => n6817, B1 => n10029, B2 => 
                           n7105, ZN => n8221);
   U9299 : AOI221_X1 port map( B1 => n9085, B2 => n10041, C1 => n9565, C2 => 
                           n10037, A => n8192, ZN => n8189);
   U9300 : OAI22_X1 port map( A1 => n10033, A2 => n6816, B1 => n10029, B2 => 
                           n7104, ZN => n8192);
   U9301 : AOI221_X1 port map( B1 => n9086, B2 => n10041, C1 => n9566, C2 => 
                           n10037, A => n8175, ZN => n8172);
   U9302 : OAI22_X1 port map( A1 => n10033, A2 => n6815, B1 => n10029, B2 => 
                           n7103, ZN => n8175);
   U9303 : AOI221_X1 port map( B1 => n9087, B2 => n10041, C1 => n9567, C2 => 
                           n10037, A => n8158, ZN => n8155);
   U9304 : OAI22_X1 port map( A1 => n10033, A2 => n6814, B1 => n10029, B2 => 
                           n7102, ZN => n8158);
   U9305 : AOI221_X1 port map( B1 => n9088, B2 => n10041, C1 => n9568, C2 => 
                           n10037, A => n8141, ZN => n8138);
   U9306 : OAI22_X1 port map( A1 => n10033, A2 => n6813, B1 => n10029, B2 => 
                           n7101, ZN => n8141);
   U9307 : AOI221_X1 port map( B1 => n9089, B2 => n10041, C1 => n9569, C2 => 
                           n10037, A => n8124, ZN => n8121);
   U9308 : OAI22_X1 port map( A1 => n10033, A2 => n6812, B1 => n10029, B2 => 
                           n7100, ZN => n8124);
   U9309 : AOI221_X1 port map( B1 => n9090, B2 => n10041, C1 => n9570, C2 => 
                           n10037, A => n8107, ZN => n8104);
   U9310 : OAI22_X1 port map( A1 => n10033, A2 => n6811, B1 => n10029, B2 => 
                           n7099, ZN => n8107);
   U9311 : AOI221_X1 port map( B1 => n9091, B2 => n10041, C1 => n9571, C2 => 
                           n10037, A => n8090, ZN => n8087);
   U9312 : OAI22_X1 port map( A1 => n10033, A2 => n6810, B1 => n10029, B2 => 
                           n7098, ZN => n8090);
   U9313 : AOI221_X1 port map( B1 => n9092, B2 => n10041, C1 => n9572, C2 => 
                           n10037, A => n8073, ZN => n8070);
   U9314 : OAI22_X1 port map( A1 => n10033, A2 => n6809, B1 => n10029, B2 => 
                           n7097, ZN => n8073);
   U9315 : AOI221_X1 port map( B1 => n9093, B2 => n10041, C1 => n9573, C2 => 
                           n10037, A => n8056, ZN => n8053);
   U9316 : OAI22_X1 port map( A1 => n10033, A2 => n6808, B1 => n10029, B2 => 
                           n7096, ZN => n8056);
   U9317 : AOI221_X1 port map( B1 => n9094, B2 => n10041, C1 => n9574, C2 => 
                           n10037, A => n8039, ZN => n8036);
   U9318 : OAI22_X1 port map( A1 => n10033, A2 => n6807, B1 => n10029, B2 => 
                           n7095, ZN => n8039);
   U9319 : AOI221_X1 port map( B1 => n9095, B2 => n10041, C1 => n9575, C2 => 
                           n10037, A => n8022, ZN => n8019);
   U9320 : OAI22_X1 port map( A1 => n10033, A2 => n6806, B1 => n10029, B2 => 
                           n7094, ZN => n8022);
   U9321 : AOI221_X1 port map( B1 => n9096, B2 => n10042, C1 => n9576, C2 => 
                           n10038, A => n8005, ZN => n8002);
   U9322 : OAI22_X1 port map( A1 => n10034, A2 => n6805, B1 => n10030, B2 => 
                           n7093, ZN => n8005);
   U9323 : AOI221_X1 port map( B1 => n9097, B2 => n10042, C1 => n9577, C2 => 
                           n10038, A => n7988, ZN => n7985);
   U9324 : OAI22_X1 port map( A1 => n10034, A2 => n6804, B1 => n10030, B2 => 
                           n7092, ZN => n7988);
   U9325 : AOI221_X1 port map( B1 => n9098, B2 => n10042, C1 => n9578, C2 => 
                           n10038, A => n7971, ZN => n7968);
   U9326 : OAI22_X1 port map( A1 => n10034, A2 => n6803, B1 => n10030, B2 => 
                           n7091, ZN => n7971);
   U9327 : AOI221_X1 port map( B1 => n9099, B2 => n10042, C1 => n9579, C2 => 
                           n10038, A => n7954, ZN => n7951);
   U9328 : OAI22_X1 port map( A1 => n10034, A2 => n6802, B1 => n10030, B2 => 
                           n7090, ZN => n7954);
   U9329 : AOI221_X1 port map( B1 => n9100, B2 => n10042, C1 => n9580, C2 => 
                           n10038, A => n7937, ZN => n7934);
   U9330 : OAI22_X1 port map( A1 => n10034, A2 => n6801, B1 => n10030, B2 => 
                           n7089, ZN => n7937);
   U9331 : AOI221_X1 port map( B1 => n9101, B2 => n10042, C1 => n9581, C2 => 
                           n10038, A => n7920, ZN => n7917);
   U9332 : OAI22_X1 port map( A1 => n10034, A2 => n6800, B1 => n10030, B2 => 
                           n7088, ZN => n7920);
   U9333 : AOI221_X1 port map( B1 => n9102, B2 => n10042, C1 => n9582, C2 => 
                           n10038, A => n7903, ZN => n7900);
   U9334 : OAI22_X1 port map( A1 => n10034, A2 => n6799, B1 => n10030, B2 => 
                           n7087, ZN => n7903);
   U9335 : AOI221_X1 port map( B1 => n9103, B2 => n10042, C1 => n9583, C2 => 
                           n10038, A => n7886, ZN => n7883);
   U9336 : OAI22_X1 port map( A1 => n10034, A2 => n6798, B1 => n10030, B2 => 
                           n7086, ZN => n7886);
   U9337 : AOI221_X1 port map( B1 => n9104, B2 => n10042, C1 => n9584, C2 => 
                           n10038, A => n7869, ZN => n7866);
   U9338 : OAI22_X1 port map( A1 => n10034, A2 => n6797, B1 => n10030, B2 => 
                           n7085, ZN => n7869);
   U9339 : AOI221_X1 port map( B1 => n9105, B2 => n10042, C1 => n9585, C2 => 
                           n10038, A => n7852, ZN => n7849);
   U9340 : OAI22_X1 port map( A1 => n10034, A2 => n6796, B1 => n10030, B2 => 
                           n7084, ZN => n7852);
   U9341 : AOI221_X1 port map( B1 => n9106, B2 => n10042, C1 => n9586, C2 => 
                           n10038, A => n7835, ZN => n7832);
   U9342 : OAI22_X1 port map( A1 => n10034, A2 => n6795, B1 => n10030, B2 => 
                           n7083, ZN => n7835);
   U9343 : AOI221_X1 port map( B1 => n9107, B2 => n10042, C1 => n9587, C2 => 
                           n10038, A => n7818, ZN => n7815);
   U9344 : OAI22_X1 port map( A1 => n10034, A2 => n6794, B1 => n10030, B2 => 
                           n7082, ZN => n7818);
   U9345 : AOI221_X1 port map( B1 => n9108, B2 => n10043, C1 => n9588, C2 => 
                           n10039, A => n7801, ZN => n7798);
   U9346 : OAI22_X1 port map( A1 => n10035, A2 => n6793, B1 => n10031, B2 => 
                           n7081, ZN => n7801);
   U9347 : AOI221_X1 port map( B1 => n9109, B2 => n10043, C1 => n9589, C2 => 
                           n10039, A => n7784, ZN => n7781);
   U9348 : OAI22_X1 port map( A1 => n10035, A2 => n6792, B1 => n10031, B2 => 
                           n7080, ZN => n7784);
   U9349 : AOI221_X1 port map( B1 => n9110, B2 => n10043, C1 => n9590, C2 => 
                           n10039, A => n7767, ZN => n7764);
   U9350 : OAI22_X1 port map( A1 => n10035, A2 => n6791, B1 => n10031, B2 => 
                           n7079, ZN => n7767);
   U9351 : AOI221_X1 port map( B1 => n9111, B2 => n10043, C1 => n9591, C2 => 
                           n10039, A => n7750, ZN => n7747);
   U9352 : OAI22_X1 port map( A1 => n10035, A2 => n6790, B1 => n10031, B2 => 
                           n7078, ZN => n7750);
   U9353 : AOI221_X1 port map( B1 => n9112, B2 => n10043, C1 => n9592, C2 => 
                           n10039, A => n7733, ZN => n7730);
   U9354 : OAI22_X1 port map( A1 => n10035, A2 => n6789, B1 => n10031, B2 => 
                           n7077, ZN => n7733);
   U9355 : AOI221_X1 port map( B1 => n9113, B2 => n10043, C1 => n9593, C2 => 
                           n10039, A => n7716, ZN => n7713);
   U9356 : OAI22_X1 port map( A1 => n10035, A2 => n6788, B1 => n10031, B2 => 
                           n7076, ZN => n7716);
   U9357 : AOI221_X1 port map( B1 => n9114, B2 => n10043, C1 => n9594, C2 => 
                           n10039, A => n7699, ZN => n7696);
   U9358 : OAI22_X1 port map( A1 => n10035, A2 => n6787, B1 => n10031, B2 => 
                           n7075, ZN => n7699);
   U9359 : AOI221_X1 port map( B1 => n9115, B2 => n10043, C1 => n9595, C2 => 
                           n10039, A => n7671, ZN => n7661);
   U9360 : OAI22_X1 port map( A1 => n10035, A2 => n6786, B1 => n10031, B2 => 
                           n7074, ZN => n7671);
   U9361 : AOI221_X1 port map( B1 => n9649, B2 => n9108, C1 => n9645, C2 => 
                           n9588, A => n8469, ZN => n8466);
   U9362 : OAI22_X1 port map( A1 => n6793, A2 => n9641, B1 => n7081, B2 => 
                           n9637, ZN => n8469);
   U9363 : AOI221_X1 port map( B1 => n9649, B2 => n9109, C1 => n9645, C2 => 
                           n9589, A => n8452, ZN => n8449);
   U9364 : OAI22_X1 port map( A1 => n6792, A2 => n9641, B1 => n7080, B2 => 
                           n9637, ZN => n8452);
   U9365 : AOI221_X1 port map( B1 => n9649, B2 => n9110, C1 => n9645, C2 => 
                           n9590, A => n8435, ZN => n8432);
   U9366 : OAI22_X1 port map( A1 => n6791, A2 => n9641, B1 => n7079, B2 => 
                           n9637, ZN => n8435);
   U9367 : AOI221_X1 port map( B1 => n9649, B2 => n9111, C1 => n9645, C2 => 
                           n9591, A => n8418, ZN => n8415);
   U9368 : OAI22_X1 port map( A1 => n6790, A2 => n9641, B1 => n7078, B2 => 
                           n9637, ZN => n8418);
   U9369 : AOI221_X1 port map( B1 => n9649, B2 => n9112, C1 => n9645, C2 => 
                           n9592, A => n8401, ZN => n8398);
   U9370 : OAI22_X1 port map( A1 => n6789, A2 => n9641, B1 => n7077, B2 => 
                           n9637, ZN => n8401);
   U9371 : AOI221_X1 port map( B1 => n9649, B2 => n9113, C1 => n9645, C2 => 
                           n9593, A => n8384, ZN => n8381);
   U9372 : OAI22_X1 port map( A1 => n6788, A2 => n9641, B1 => n7076, B2 => 
                           n9637, ZN => n8384);
   U9373 : AOI221_X1 port map( B1 => n9649, B2 => n9114, C1 => n9645, C2 => 
                           n9594, A => n8367, ZN => n8364);
   U9374 : OAI22_X1 port map( A1 => n6787, A2 => n9641, B1 => n7075, B2 => 
                           n9637, ZN => n8367);
   U9375 : AOI221_X1 port map( B1 => n9649, B2 => n9115, C1 => n9645, C2 => 
                           n9595, A => n8339, ZN => n8329);
   U9376 : OAI22_X1 port map( A1 => n6786, A2 => n9641, B1 => n7074, B2 => 
                           n9637, ZN => n8339);
   U9377 : AOI221_X1 port map( B1 => n9647, B2 => n9084, C1 => n9643, C2 => 
                           n9564, A => n8889, ZN => n8884);
   U9378 : OAI22_X1 port map( A1 => n6817, A2 => n9639, B1 => n7105, B2 => 
                           n9635, ZN => n8889);
   U9379 : AOI221_X1 port map( B1 => n9647, B2 => n9085, C1 => n9643, C2 => 
                           n9565, A => n8860, ZN => n8857);
   U9380 : OAI22_X1 port map( A1 => n6816, A2 => n9639, B1 => n7104, B2 => 
                           n9635, ZN => n8860);
   U9381 : AOI221_X1 port map( B1 => n9647, B2 => n9086, C1 => n9643, C2 => 
                           n9566, A => n8843, ZN => n8840);
   U9382 : OAI22_X1 port map( A1 => n6815, A2 => n9639, B1 => n7103, B2 => 
                           n9635, ZN => n8843);
   U9383 : AOI221_X1 port map( B1 => n9647, B2 => n9087, C1 => n9643, C2 => 
                           n9567, A => n8826, ZN => n8823);
   U9384 : OAI22_X1 port map( A1 => n6814, A2 => n9639, B1 => n7102, B2 => 
                           n9635, ZN => n8826);
   U9385 : AOI221_X1 port map( B1 => n9647, B2 => n9088, C1 => n9643, C2 => 
                           n9568, A => n8809, ZN => n8806);
   U9386 : OAI22_X1 port map( A1 => n6813, A2 => n9639, B1 => n7101, B2 => 
                           n9635, ZN => n8809);
   U9387 : AOI221_X1 port map( B1 => n9647, B2 => n9089, C1 => n9643, C2 => 
                           n9569, A => n8792, ZN => n8789);
   U9388 : OAI22_X1 port map( A1 => n6812, A2 => n9639, B1 => n7100, B2 => 
                           n9635, ZN => n8792);
   U9389 : AOI221_X1 port map( B1 => n9647, B2 => n9090, C1 => n9643, C2 => 
                           n9570, A => n8775, ZN => n8772);
   U9390 : OAI22_X1 port map( A1 => n6811, A2 => n9639, B1 => n7099, B2 => 
                           n9635, ZN => n8775);
   U9391 : AOI221_X1 port map( B1 => n9647, B2 => n9091, C1 => n9643, C2 => 
                           n9571, A => n8758, ZN => n8755);
   U9392 : OAI22_X1 port map( A1 => n6810, A2 => n9639, B1 => n7098, B2 => 
                           n9635, ZN => n8758);
   U9393 : AOI221_X1 port map( B1 => n9647, B2 => n9092, C1 => n9643, C2 => 
                           n9572, A => n8741, ZN => n8738);
   U9394 : OAI22_X1 port map( A1 => n6809, A2 => n9639, B1 => n7097, B2 => 
                           n9635, ZN => n8741);
   U9395 : AOI221_X1 port map( B1 => n9647, B2 => n9093, C1 => n9643, C2 => 
                           n9573, A => n8724, ZN => n8721);
   U9396 : OAI22_X1 port map( A1 => n6808, A2 => n9639, B1 => n7096, B2 => 
                           n9635, ZN => n8724);
   U9397 : AOI221_X1 port map( B1 => n9647, B2 => n9094, C1 => n9643, C2 => 
                           n9574, A => n8707, ZN => n8704);
   U9398 : OAI22_X1 port map( A1 => n6807, A2 => n9639, B1 => n7095, B2 => 
                           n9635, ZN => n8707);
   U9399 : AOI221_X1 port map( B1 => n9647, B2 => n9095, C1 => n9643, C2 => 
                           n9575, A => n8690, ZN => n8687);
   U9400 : OAI22_X1 port map( A1 => n6806, A2 => n9639, B1 => n7094, B2 => 
                           n9635, ZN => n8690);
   U9401 : AOI221_X1 port map( B1 => n9648, B2 => n9096, C1 => n9644, C2 => 
                           n9576, A => n8673, ZN => n8670);
   U9402 : OAI22_X1 port map( A1 => n6805, A2 => n9640, B1 => n7093, B2 => 
                           n9636, ZN => n8673);
   U9403 : AOI221_X1 port map( B1 => n9648, B2 => n9097, C1 => n9644, C2 => 
                           n9577, A => n8656, ZN => n8653);
   U9404 : OAI22_X1 port map( A1 => n6804, A2 => n9640, B1 => n7092, B2 => 
                           n9636, ZN => n8656);
   U9405 : AOI221_X1 port map( B1 => n9648, B2 => n9098, C1 => n9644, C2 => 
                           n9578, A => n8639, ZN => n8636);
   U9406 : OAI22_X1 port map( A1 => n6803, A2 => n9640, B1 => n7091, B2 => 
                           n9636, ZN => n8639);
   U9407 : AOI221_X1 port map( B1 => n9648, B2 => n9099, C1 => n9644, C2 => 
                           n9579, A => n8622, ZN => n8619);
   U9408 : OAI22_X1 port map( A1 => n6802, A2 => n9640, B1 => n7090, B2 => 
                           n9636, ZN => n8622);
   U9409 : AOI221_X1 port map( B1 => n9648, B2 => n9100, C1 => n9644, C2 => 
                           n9580, A => n8605, ZN => n8602);
   U9410 : OAI22_X1 port map( A1 => n6801, A2 => n9640, B1 => n7089, B2 => 
                           n9636, ZN => n8605);
   U9411 : AOI221_X1 port map( B1 => n9648, B2 => n9101, C1 => n9644, C2 => 
                           n9581, A => n8588, ZN => n8585);
   U9412 : OAI22_X1 port map( A1 => n6800, A2 => n9640, B1 => n7088, B2 => 
                           n9636, ZN => n8588);
   U9413 : AOI221_X1 port map( B1 => n9648, B2 => n9102, C1 => n9644, C2 => 
                           n9582, A => n8571, ZN => n8568);
   U9414 : OAI22_X1 port map( A1 => n6799, A2 => n9640, B1 => n7087, B2 => 
                           n9636, ZN => n8571);
   U9415 : AOI221_X1 port map( B1 => n9648, B2 => n9103, C1 => n9644, C2 => 
                           n9583, A => n8554, ZN => n8551);
   U9416 : OAI22_X1 port map( A1 => n6798, A2 => n9640, B1 => n7086, B2 => 
                           n9636, ZN => n8554);
   U9417 : AOI221_X1 port map( B1 => n9648, B2 => n9104, C1 => n9644, C2 => 
                           n9584, A => n8537, ZN => n8534);
   U9418 : OAI22_X1 port map( A1 => n6797, A2 => n9640, B1 => n7085, B2 => 
                           n9636, ZN => n8537);
   U9419 : AOI221_X1 port map( B1 => n9648, B2 => n9105, C1 => n9644, C2 => 
                           n9585, A => n8520, ZN => n8517);
   U9420 : OAI22_X1 port map( A1 => n6796, A2 => n9640, B1 => n7084, B2 => 
                           n9636, ZN => n8520);
   U9421 : AOI221_X1 port map( B1 => n9648, B2 => n9106, C1 => n9644, C2 => 
                           n9586, A => n8503, ZN => n8500);
   U9422 : OAI22_X1 port map( A1 => n6795, A2 => n9640, B1 => n7083, B2 => 
                           n9636, ZN => n8503);
   U9423 : AOI221_X1 port map( B1 => n9648, B2 => n9107, C1 => n9644, C2 => 
                           n9587, A => n8486, ZN => n8483);
   U9424 : OAI22_X1 port map( A1 => n6794, A2 => n9640, B1 => n7082, B2 => 
                           n9636, ZN => n8486);
   U9425 : OAI22_X1 port map( A1 => n480, A2 => n9603, B1 => n544, B2 => n9599,
                           ZN => n8891);
   U9426 : OAI22_X1 port map( A1 => n481, A2 => n9603, B1 => n545, B2 => n9599,
                           ZN => n8862);
   U9427 : OAI22_X1 port map( A1 => n482, A2 => n9603, B1 => n546, B2 => n9599,
                           ZN => n8845);
   U9428 : OAI22_X1 port map( A1 => n483, A2 => n9603, B1 => n547, B2 => n9599,
                           ZN => n8828);
   U9429 : OAI22_X1 port map( A1 => n484, A2 => n9603, B1 => n548, B2 => n9599,
                           ZN => n8811);
   U9430 : OAI22_X1 port map( A1 => n485, A2 => n9603, B1 => n549, B2 => n9599,
                           ZN => n8794);
   U9431 : OAI22_X1 port map( A1 => n486, A2 => n9603, B1 => n550, B2 => n9599,
                           ZN => n8777);
   U9432 : OAI22_X1 port map( A1 => n487, A2 => n9603, B1 => n551, B2 => n9599,
                           ZN => n8760);
   U9433 : OAI22_X1 port map( A1 => n488, A2 => n9603, B1 => n552, B2 => n9599,
                           ZN => n8743);
   U9434 : OAI22_X1 port map( A1 => n489, A2 => n9603, B1 => n553, B2 => n9599,
                           ZN => n8726);
   U9435 : OAI22_X1 port map( A1 => n490, A2 => n9603, B1 => n554, B2 => n9599,
                           ZN => n8709);
   U9436 : OAI22_X1 port map( A1 => n491, A2 => n9603, B1 => n555, B2 => n9599,
                           ZN => n8692);
   U9437 : OAI22_X1 port map( A1 => n492, A2 => n9604, B1 => n556, B2 => n9600,
                           ZN => n8675);
   U9438 : OAI22_X1 port map( A1 => n493, A2 => n9604, B1 => n557, B2 => n9600,
                           ZN => n8658);
   U9439 : OAI22_X1 port map( A1 => n494, A2 => n9604, B1 => n558, B2 => n9600,
                           ZN => n8641);
   U9440 : OAI22_X1 port map( A1 => n495, A2 => n9604, B1 => n559, B2 => n9600,
                           ZN => n8624);
   U9441 : OAI22_X1 port map( A1 => n496, A2 => n9604, B1 => n560, B2 => n9600,
                           ZN => n8607);
   U9442 : OAI22_X1 port map( A1 => n497, A2 => n9604, B1 => n561, B2 => n9600,
                           ZN => n8590);
   U9443 : OAI22_X1 port map( A1 => n498, A2 => n9604, B1 => n562, B2 => n9600,
                           ZN => n8573);
   U9444 : OAI22_X1 port map( A1 => n499, A2 => n9604, B1 => n563, B2 => n9600,
                           ZN => n8556);
   U9445 : OAI22_X1 port map( A1 => n500, A2 => n9604, B1 => n564, B2 => n9600,
                           ZN => n8539);
   U9446 : OAI22_X1 port map( A1 => n501, A2 => n9604, B1 => n565, B2 => n9600,
                           ZN => n8522);
   U9447 : OAI22_X1 port map( A1 => n502, A2 => n9604, B1 => n566, B2 => n9600,
                           ZN => n8505);
   U9448 : OAI22_X1 port map( A1 => n503, A2 => n9604, B1 => n567, B2 => n9600,
                           ZN => n8488);
   U9449 : OAI22_X1 port map( A1 => n504, A2 => n9605, B1 => n568, B2 => n9601,
                           ZN => n8471);
   U9450 : OAI22_X1 port map( A1 => n505, A2 => n9605, B1 => n569, B2 => n9601,
                           ZN => n8454);
   U9451 : OAI22_X1 port map( A1 => n506, A2 => n9605, B1 => n570, B2 => n9601,
                           ZN => n8437);
   U9452 : OAI22_X1 port map( A1 => n507, A2 => n9605, B1 => n571, B2 => n9601,
                           ZN => n8420);
   U9453 : OAI22_X1 port map( A1 => n508, A2 => n9605, B1 => n572, B2 => n9601,
                           ZN => n8403);
   U9454 : OAI22_X1 port map( A1 => n509, A2 => n9605, B1 => n573, B2 => n9601,
                           ZN => n8386);
   U9455 : OAI22_X1 port map( A1 => n510, A2 => n9605, B1 => n574, B2 => n9601,
                           ZN => n8369);
   U9456 : OAI22_X1 port map( A1 => n511, A2 => n9605, B1 => n575, B2 => n9601,
                           ZN => n8350);
   U9457 : OAI22_X1 port map( A1 => n480, A2 => n9997, B1 => n544, B2 => n9993,
                           ZN => n8223);
   U9458 : OAI22_X1 port map( A1 => n481, A2 => n9997, B1 => n545, B2 => n9993,
                           ZN => n8194);
   U9459 : OAI22_X1 port map( A1 => n482, A2 => n9997, B1 => n546, B2 => n9993,
                           ZN => n8177);
   U9460 : OAI22_X1 port map( A1 => n483, A2 => n9997, B1 => n547, B2 => n9993,
                           ZN => n8160);
   U9461 : OAI22_X1 port map( A1 => n484, A2 => n9997, B1 => n548, B2 => n9993,
                           ZN => n8143);
   U9462 : OAI22_X1 port map( A1 => n485, A2 => n9997, B1 => n549, B2 => n9993,
                           ZN => n8126);
   U9463 : OAI22_X1 port map( A1 => n486, A2 => n9997, B1 => n550, B2 => n9993,
                           ZN => n8109);
   U9464 : OAI22_X1 port map( A1 => n487, A2 => n9997, B1 => n551, B2 => n9993,
                           ZN => n8092);
   U9465 : OAI22_X1 port map( A1 => n488, A2 => n9997, B1 => n552, B2 => n9993,
                           ZN => n8075);
   U9466 : OAI22_X1 port map( A1 => n489, A2 => n9997, B1 => n553, B2 => n9993,
                           ZN => n8058);
   U9467 : OAI22_X1 port map( A1 => n490, A2 => n9997, B1 => n554, B2 => n9993,
                           ZN => n8041);
   U9468 : OAI22_X1 port map( A1 => n491, A2 => n9997, B1 => n555, B2 => n9993,
                           ZN => n8024);
   U9469 : OAI22_X1 port map( A1 => n492, A2 => n9998, B1 => n556, B2 => n9994,
                           ZN => n8007);
   U9470 : OAI22_X1 port map( A1 => n493, A2 => n9998, B1 => n557, B2 => n9994,
                           ZN => n7990);
   U9471 : OAI22_X1 port map( A1 => n494, A2 => n9998, B1 => n558, B2 => n9994,
                           ZN => n7973);
   U9472 : OAI22_X1 port map( A1 => n495, A2 => n9998, B1 => n559, B2 => n9994,
                           ZN => n7956);
   U9473 : OAI22_X1 port map( A1 => n496, A2 => n9998, B1 => n560, B2 => n9994,
                           ZN => n7939);
   U9474 : OAI22_X1 port map( A1 => n497, A2 => n9998, B1 => n561, B2 => n9994,
                           ZN => n7922);
   U9475 : OAI22_X1 port map( A1 => n498, A2 => n9998, B1 => n562, B2 => n9994,
                           ZN => n7905);
   U9476 : OAI22_X1 port map( A1 => n499, A2 => n9998, B1 => n563, B2 => n9994,
                           ZN => n7888);
   U9477 : OAI22_X1 port map( A1 => n500, A2 => n9998, B1 => n564, B2 => n9994,
                           ZN => n7871);
   U9478 : OAI22_X1 port map( A1 => n501, A2 => n9998, B1 => n565, B2 => n9994,
                           ZN => n7854);
   U9479 : OAI22_X1 port map( A1 => n502, A2 => n9998, B1 => n566, B2 => n9994,
                           ZN => n7837);
   U9480 : OAI22_X1 port map( A1 => n503, A2 => n9998, B1 => n567, B2 => n9994,
                           ZN => n7820);
   U9481 : OAI22_X1 port map( A1 => n504, A2 => n9999, B1 => n568, B2 => n9995,
                           ZN => n7803);
   U9482 : OAI22_X1 port map( A1 => n505, A2 => n9999, B1 => n569, B2 => n9995,
                           ZN => n7786);
   U9483 : OAI22_X1 port map( A1 => n506, A2 => n9999, B1 => n570, B2 => n9995,
                           ZN => n7769);
   U9484 : OAI22_X1 port map( A1 => n507, A2 => n9999, B1 => n571, B2 => n9995,
                           ZN => n7752);
   U9485 : OAI22_X1 port map( A1 => n508, A2 => n9999, B1 => n572, B2 => n9995,
                           ZN => n7735);
   U9486 : OAI22_X1 port map( A1 => n509, A2 => n9999, B1 => n573, B2 => n9995,
                           ZN => n7718);
   U9487 : OAI22_X1 port map( A1 => n510, A2 => n9999, B1 => n574, B2 => n9995,
                           ZN => n7701);
   U9488 : OAI22_X1 port map( A1 => n511, A2 => n9999, B1 => n575, B2 => n9995,
                           ZN => n7682);
   U9489 : OAI22_X1 port map( A1 => n640, A2 => n10102, B1 => n10098, B2 => 
                           n7360, ZN => n8205);
   U9490 : OAI22_X1 port map( A1 => n641, A2 => n10102, B1 => n10098, B2 => 
                           n7359, ZN => n8183);
   U9491 : OAI22_X1 port map( A1 => n642, A2 => n10102, B1 => n10098, B2 => 
                           n7358, ZN => n8166);
   U9492 : OAI22_X1 port map( A1 => n643, A2 => n10102, B1 => n10098, B2 => 
                           n7357, ZN => n8149);
   U9493 : OAI22_X1 port map( A1 => n644, A2 => n10102, B1 => n10098, B2 => 
                           n7356, ZN => n8132);
   U9494 : OAI22_X1 port map( A1 => n645, A2 => n10102, B1 => n10098, B2 => 
                           n7355, ZN => n8115);
   U9495 : OAI22_X1 port map( A1 => n646, A2 => n10102, B1 => n10098, B2 => 
                           n7354, ZN => n8098);
   U9496 : OAI22_X1 port map( A1 => n647, A2 => n10102, B1 => n10098, B2 => 
                           n7353, ZN => n8081);
   U9497 : OAI22_X1 port map( A1 => n648, A2 => n10102, B1 => n10098, B2 => 
                           n7352, ZN => n8064);
   U9498 : OAI22_X1 port map( A1 => n649, A2 => n10102, B1 => n10098, B2 => 
                           n7351, ZN => n8047);
   U9499 : OAI22_X1 port map( A1 => n650, A2 => n10102, B1 => n10098, B2 => 
                           n7350, ZN => n8030);
   U9500 : OAI22_X1 port map( A1 => n651, A2 => n10102, B1 => n10098, B2 => 
                           n7349, ZN => n8013);
   U9501 : OAI22_X1 port map( A1 => n652, A2 => n10103, B1 => n10099, B2 => 
                           n7348, ZN => n7996);
   U9502 : OAI22_X1 port map( A1 => n653, A2 => n10103, B1 => n10099, B2 => 
                           n7347, ZN => n7979);
   U9503 : OAI22_X1 port map( A1 => n654, A2 => n10103, B1 => n10099, B2 => 
                           n7346, ZN => n7962);
   U9504 : OAI22_X1 port map( A1 => n655, A2 => n10103, B1 => n10099, B2 => 
                           n7345, ZN => n7945);
   U9505 : OAI22_X1 port map( A1 => n656, A2 => n10103, B1 => n10099, B2 => 
                           n7344, ZN => n7928);
   U9506 : OAI22_X1 port map( A1 => n657, A2 => n10103, B1 => n10099, B2 => 
                           n7343, ZN => n7911);
   U9507 : OAI22_X1 port map( A1 => n658, A2 => n10103, B1 => n10099, B2 => 
                           n7342, ZN => n7894);
   U9508 : OAI22_X1 port map( A1 => n659, A2 => n10103, B1 => n10099, B2 => 
                           n7341, ZN => n7877);
   U9509 : OAI22_X1 port map( A1 => n660, A2 => n10103, B1 => n10099, B2 => 
                           n7340, ZN => n7860);
   U9510 : OAI22_X1 port map( A1 => n661, A2 => n10103, B1 => n10099, B2 => 
                           n7339, ZN => n7843);
   U9511 : OAI22_X1 port map( A1 => n662, A2 => n10103, B1 => n10099, B2 => 
                           n7338, ZN => n7826);
   U9512 : OAI22_X1 port map( A1 => n663, A2 => n10103, B1 => n10099, B2 => 
                           n7337, ZN => n7809);
   U9513 : OAI22_X1 port map( A1 => n664, A2 => n10104, B1 => n10100, B2 => 
                           n7336, ZN => n7792);
   U9514 : OAI22_X1 port map( A1 => n665, A2 => n10104, B1 => n10100, B2 => 
                           n7335, ZN => n7775);
   U9515 : OAI22_X1 port map( A1 => n666, A2 => n10104, B1 => n10100, B2 => 
                           n7334, ZN => n7758);
   U9516 : OAI22_X1 port map( A1 => n667, A2 => n10104, B1 => n10100, B2 => 
                           n7333, ZN => n7741);
   U9517 : OAI22_X1 port map( A1 => n668, A2 => n10104, B1 => n10100, B2 => 
                           n7332, ZN => n7724);
   U9518 : OAI22_X1 port map( A1 => n669, A2 => n10104, B1 => n10100, B2 => 
                           n7331, ZN => n7707);
   U9519 : OAI22_X1 port map( A1 => n670, A2 => n10104, B1 => n10100, B2 => 
                           n7330, ZN => n7690);
   U9520 : OAI22_X1 port map( A1 => n671, A2 => n10104, B1 => n10100, B2 => 
                           n7329, ZN => n7645);
   U9521 : OAI22_X1 port map( A1 => n464, A2 => n10087, B1 => n10083, B2 => 
                           n7376, ZN => n7929);
   U9522 : OAI22_X1 port map( A1 => n465, A2 => n10087, B1 => n10083, B2 => 
                           n7375, ZN => n7912);
   U9523 : OAI22_X1 port map( A1 => n466, A2 => n10087, B1 => n10083, B2 => 
                           n7374, ZN => n7895);
   U9524 : OAI22_X1 port map( A1 => n467, A2 => n10087, B1 => n10083, B2 => 
                           n7373, ZN => n7878);
   U9525 : OAI22_X1 port map( A1 => n468, A2 => n10086, B1 => n10083, B2 => 
                           n7372, ZN => n7861);
   U9526 : OAI22_X1 port map( A1 => n469, A2 => n10086, B1 => n10083, B2 => 
                           n7371, ZN => n7844);
   U9527 : OAI22_X1 port map( A1 => n470, A2 => n10086, B1 => n10083, B2 => 
                           n7370, ZN => n7827);
   U9528 : OAI22_X1 port map( A1 => n471, A2 => n10086, B1 => n10083, B2 => 
                           n7369, ZN => n7810);
   U9529 : OAI22_X1 port map( A1 => n472, A2 => n10086, B1 => n10084, B2 => 
                           n7368, ZN => n7793);
   U9530 : OAI22_X1 port map( A1 => n473, A2 => n10086, B1 => n10084, B2 => 
                           n7367, ZN => n7776);
   U9531 : OAI22_X1 port map( A1 => n474, A2 => n10086, B1 => n10084, B2 => 
                           n7366, ZN => n7759);
   U9532 : OAI22_X1 port map( A1 => n475, A2 => n10086, B1 => n10084, B2 => 
                           n7365, ZN => n7742);
   U9533 : OAI22_X1 port map( A1 => n476, A2 => n10086, B1 => n10084, B2 => 
                           n7364, ZN => n7725);
   U9534 : OAI22_X1 port map( A1 => n477, A2 => n10086, B1 => n10084, B2 => 
                           n7363, ZN => n7708);
   U9535 : OAI22_X1 port map( A1 => n478, A2 => n10086, B1 => n10084, B2 => 
                           n7362, ZN => n7691);
   U9536 : OAI22_X1 port map( A1 => n479, A2 => n10086, B1 => n10084, B2 => 
                           n7361, ZN => n7650);
   U9537 : OAI22_X1 port map( A1 => n640, A2 => n9708, B1 => n7360, B2 => n9704
                           , ZN => n8873);
   U9538 : OAI22_X1 port map( A1 => n641, A2 => n9708, B1 => n7359, B2 => n9704
                           , ZN => n8851);
   U9539 : OAI22_X1 port map( A1 => n642, A2 => n9708, B1 => n7358, B2 => n9704
                           , ZN => n8834);
   U9540 : OAI22_X1 port map( A1 => n643, A2 => n9708, B1 => n7357, B2 => n9704
                           , ZN => n8817);
   U9541 : OAI22_X1 port map( A1 => n644, A2 => n9708, B1 => n7356, B2 => n9704
                           , ZN => n8800);
   U9542 : OAI22_X1 port map( A1 => n645, A2 => n9708, B1 => n7355, B2 => n9704
                           , ZN => n8783);
   U9543 : OAI22_X1 port map( A1 => n646, A2 => n9708, B1 => n7354, B2 => n9704
                           , ZN => n8766);
   U9544 : OAI22_X1 port map( A1 => n647, A2 => n9708, B1 => n7353, B2 => n9704
                           , ZN => n8749);
   U9545 : OAI22_X1 port map( A1 => n648, A2 => n9708, B1 => n7352, B2 => n9704
                           , ZN => n8732);
   U9546 : OAI22_X1 port map( A1 => n649, A2 => n9708, B1 => n7351, B2 => n9704
                           , ZN => n8715);
   U9547 : OAI22_X1 port map( A1 => n650, A2 => n9708, B1 => n7350, B2 => n9704
                           , ZN => n8698);
   U9548 : OAI22_X1 port map( A1 => n651, A2 => n9708, B1 => n7349, B2 => n9704
                           , ZN => n8681);
   U9549 : OAI22_X1 port map( A1 => n652, A2 => n9709, B1 => n7348, B2 => n9705
                           , ZN => n8664);
   U9550 : OAI22_X1 port map( A1 => n653, A2 => n9709, B1 => n7347, B2 => n9705
                           , ZN => n8647);
   U9551 : OAI22_X1 port map( A1 => n654, A2 => n9709, B1 => n7346, B2 => n9705
                           , ZN => n8630);
   U9552 : OAI22_X1 port map( A1 => n655, A2 => n9709, B1 => n7345, B2 => n9705
                           , ZN => n8613);
   U9553 : OAI22_X1 port map( A1 => n656, A2 => n9709, B1 => n7344, B2 => n9705
                           , ZN => n8596);
   U9554 : OAI22_X1 port map( A1 => n657, A2 => n9709, B1 => n7343, B2 => n9705
                           , ZN => n8579);
   U9555 : OAI22_X1 port map( A1 => n658, A2 => n9709, B1 => n7342, B2 => n9705
                           , ZN => n8562);
   U9556 : OAI22_X1 port map( A1 => n659, A2 => n9709, B1 => n7341, B2 => n9705
                           , ZN => n8545);
   U9557 : OAI22_X1 port map( A1 => n660, A2 => n9709, B1 => n7340, B2 => n9705
                           , ZN => n8528);
   U9558 : OAI22_X1 port map( A1 => n661, A2 => n9709, B1 => n7339, B2 => n9705
                           , ZN => n8511);
   U9559 : OAI22_X1 port map( A1 => n662, A2 => n9709, B1 => n7338, B2 => n9705
                           , ZN => n8494);
   U9560 : OAI22_X1 port map( A1 => n663, A2 => n9709, B1 => n7337, B2 => n9705
                           , ZN => n8477);
   U9561 : OAI22_X1 port map( A1 => n664, A2 => n9710, B1 => n7336, B2 => n9706
                           , ZN => n8460);
   U9562 : OAI22_X1 port map( A1 => n665, A2 => n9710, B1 => n7335, B2 => n9706
                           , ZN => n8443);
   U9563 : OAI22_X1 port map( A1 => n666, A2 => n9710, B1 => n7334, B2 => n9706
                           , ZN => n8426);
   U9564 : OAI22_X1 port map( A1 => n667, A2 => n9710, B1 => n7333, B2 => n9706
                           , ZN => n8409);
   U9565 : OAI22_X1 port map( A1 => n668, A2 => n9710, B1 => n7332, B2 => n9706
                           , ZN => n8392);
   U9566 : OAI22_X1 port map( A1 => n669, A2 => n9710, B1 => n7331, B2 => n9706
                           , ZN => n8375);
   U9567 : OAI22_X1 port map( A1 => n670, A2 => n9710, B1 => n7330, B2 => n9706
                           , ZN => n8358);
   U9568 : OAI22_X1 port map( A1 => n671, A2 => n9710, B1 => n7329, B2 => n9706
                           , ZN => n8313);
   U9569 : OAI22_X1 port map( A1 => n464, A2 => n9693, B1 => n7376, B2 => n9689
                           , ZN => n8597);
   U9570 : OAI22_X1 port map( A1 => n465, A2 => n9693, B1 => n7375, B2 => n9689
                           , ZN => n8580);
   U9571 : OAI22_X1 port map( A1 => n466, A2 => n9693, B1 => n7374, B2 => n9689
                           , ZN => n8563);
   U9572 : OAI22_X1 port map( A1 => n467, A2 => n9693, B1 => n7373, B2 => n9689
                           , ZN => n8546);
   U9573 : OAI22_X1 port map( A1 => n468, A2 => n9693, B1 => n7372, B2 => n9689
                           , ZN => n8529);
   U9574 : OAI22_X1 port map( A1 => n469, A2 => n9693, B1 => n7371, B2 => n9689
                           , ZN => n8512);
   U9575 : OAI22_X1 port map( A1 => n470, A2 => n9693, B1 => n7370, B2 => n9689
                           , ZN => n8495);
   U9576 : OAI22_X1 port map( A1 => n471, A2 => n9693, B1 => n7369, B2 => n9689
                           , ZN => n8478);
   U9577 : OAI22_X1 port map( A1 => n472, A2 => n9694, B1 => n7368, B2 => n9690
                           , ZN => n8461);
   U9578 : OAI22_X1 port map( A1 => n473, A2 => n9694, B1 => n7367, B2 => n9690
                           , ZN => n8444);
   U9579 : OAI22_X1 port map( A1 => n474, A2 => n9694, B1 => n7366, B2 => n9690
                           , ZN => n8427);
   U9580 : OAI22_X1 port map( A1 => n475, A2 => n9694, B1 => n7365, B2 => n9690
                           , ZN => n8410);
   U9581 : OAI22_X1 port map( A1 => n476, A2 => n9694, B1 => n7364, B2 => n9690
                           , ZN => n8393);
   U9582 : OAI22_X1 port map( A1 => n477, A2 => n9694, B1 => n7363, B2 => n9690
                           , ZN => n8376);
   U9583 : OAI22_X1 port map( A1 => n478, A2 => n9694, B1 => n7362, B2 => n9690
                           , ZN => n8359);
   U9584 : OAI22_X1 port map( A1 => n479, A2 => n9694, B1 => n7361, B2 => n9690
                           , ZN => n8318);
   U9585 : OAI22_X1 port map( A1 => n704, A2 => n9724, B1 => n512, B2 => n9720,
                           ZN => n8867);
   U9586 : OAI22_X1 port map( A1 => n705, A2 => n9724, B1 => n513, B2 => n9720,
                           ZN => n8850);
   U9587 : OAI22_X1 port map( A1 => n706, A2 => n9724, B1 => n514, B2 => n9720,
                           ZN => n8833);
   U9588 : OAI22_X1 port map( A1 => n707, A2 => n9724, B1 => n515, B2 => n9720,
                           ZN => n8816);
   U9589 : OAI22_X1 port map( A1 => n708, A2 => n9724, B1 => n516, B2 => n9720,
                           ZN => n8799);
   U9590 : OAI22_X1 port map( A1 => n709, A2 => n9724, B1 => n517, B2 => n9720,
                           ZN => n8782);
   U9591 : OAI22_X1 port map( A1 => n710, A2 => n9724, B1 => n518, B2 => n9720,
                           ZN => n8765);
   U9592 : OAI22_X1 port map( A1 => n711, A2 => n9724, B1 => n519, B2 => n9720,
                           ZN => n8748);
   U9593 : OAI22_X1 port map( A1 => n712, A2 => n9724, B1 => n520, B2 => n9720,
                           ZN => n8731);
   U9594 : OAI22_X1 port map( A1 => n713, A2 => n9724, B1 => n521, B2 => n9720,
                           ZN => n8714);
   U9595 : OAI22_X1 port map( A1 => n714, A2 => n9724, B1 => n522, B2 => n9720,
                           ZN => n8697);
   U9596 : OAI22_X1 port map( A1 => n715, A2 => n9724, B1 => n523, B2 => n9720,
                           ZN => n8680);
   U9597 : OAI22_X1 port map( A1 => n716, A2 => n9725, B1 => n524, B2 => n9721,
                           ZN => n8663);
   U9598 : OAI22_X1 port map( A1 => n717, A2 => n9725, B1 => n525, B2 => n9721,
                           ZN => n8646);
   U9599 : OAI22_X1 port map( A1 => n718, A2 => n9725, B1 => n526, B2 => n9721,
                           ZN => n8629);
   U9600 : OAI22_X1 port map( A1 => n719, A2 => n9725, B1 => n527, B2 => n9721,
                           ZN => n8612);
   U9601 : OAI22_X1 port map( A1 => n720, A2 => n9725, B1 => n528, B2 => n9721,
                           ZN => n8595);
   U9602 : OAI22_X1 port map( A1 => n721, A2 => n9725, B1 => n529, B2 => n9721,
                           ZN => n8578);
   U9603 : OAI22_X1 port map( A1 => n722, A2 => n9725, B1 => n530, B2 => n9721,
                           ZN => n8561);
   U9604 : OAI22_X1 port map( A1 => n723, A2 => n9725, B1 => n531, B2 => n9721,
                           ZN => n8544);
   U9605 : OAI22_X1 port map( A1 => n724, A2 => n9725, B1 => n532, B2 => n9721,
                           ZN => n8527);
   U9606 : OAI22_X1 port map( A1 => n725, A2 => n9725, B1 => n533, B2 => n9721,
                           ZN => n8510);
   U9607 : OAI22_X1 port map( A1 => n726, A2 => n9725, B1 => n534, B2 => n9721,
                           ZN => n8493);
   U9608 : OAI22_X1 port map( A1 => n727, A2 => n9725, B1 => n535, B2 => n9721,
                           ZN => n8476);
   U9609 : OAI22_X1 port map( A1 => n728, A2 => n9726, B1 => n536, B2 => n9722,
                           ZN => n8459);
   U9610 : OAI22_X1 port map( A1 => n729, A2 => n9726, B1 => n537, B2 => n9722,
                           ZN => n8442);
   U9611 : OAI22_X1 port map( A1 => n730, A2 => n9726, B1 => n538, B2 => n9722,
                           ZN => n8425);
   U9612 : OAI22_X1 port map( A1 => n731, A2 => n9726, B1 => n539, B2 => n9722,
                           ZN => n8408);
   U9613 : OAI22_X1 port map( A1 => n732, A2 => n9726, B1 => n540, B2 => n9722,
                           ZN => n8391);
   U9614 : OAI22_X1 port map( A1 => n733, A2 => n9726, B1 => n541, B2 => n9722,
                           ZN => n8374);
   U9615 : OAI22_X1 port map( A1 => n734, A2 => n9726, B1 => n542, B2 => n9722,
                           ZN => n8357);
   U9616 : OAI22_X1 port map( A1 => n735, A2 => n9726, B1 => n543, B2 => n9722,
                           ZN => n8308);
   U9617 : OAI22_X1 port map( A1 => n704, A2 => n10118, B1 => n512, B2 => 
                           n10114, ZN => n8199);
   U9618 : OAI22_X1 port map( A1 => n705, A2 => n10118, B1 => n513, B2 => 
                           n10114, ZN => n8182);
   U9619 : OAI22_X1 port map( A1 => n706, A2 => n10118, B1 => n514, B2 => 
                           n10114, ZN => n8165);
   U9620 : OAI22_X1 port map( A1 => n707, A2 => n10118, B1 => n515, B2 => 
                           n10114, ZN => n8148);
   U9621 : OAI22_X1 port map( A1 => n708, A2 => n10118, B1 => n516, B2 => 
                           n10114, ZN => n8131);
   U9622 : OAI22_X1 port map( A1 => n709, A2 => n10118, B1 => n517, B2 => 
                           n10114, ZN => n8114);
   U9623 : OAI22_X1 port map( A1 => n710, A2 => n10118, B1 => n518, B2 => 
                           n10114, ZN => n8097);
   U9624 : OAI22_X1 port map( A1 => n711, A2 => n10118, B1 => n519, B2 => 
                           n10114, ZN => n8080);
   U9625 : OAI22_X1 port map( A1 => n712, A2 => n10118, B1 => n520, B2 => 
                           n10114, ZN => n8063);
   U9626 : OAI22_X1 port map( A1 => n713, A2 => n10118, B1 => n521, B2 => 
                           n10114, ZN => n8046);
   U9627 : OAI22_X1 port map( A1 => n714, A2 => n10118, B1 => n522, B2 => 
                           n10114, ZN => n8029);
   U9628 : OAI22_X1 port map( A1 => n715, A2 => n10118, B1 => n523, B2 => 
                           n10114, ZN => n8012);
   U9629 : OAI22_X1 port map( A1 => n716, A2 => n10119, B1 => n524, B2 => 
                           n10115, ZN => n7995);
   U9630 : OAI22_X1 port map( A1 => n717, A2 => n10119, B1 => n525, B2 => 
                           n10115, ZN => n7978);
   U9631 : OAI22_X1 port map( A1 => n718, A2 => n10119, B1 => n526, B2 => 
                           n10115, ZN => n7961);
   U9632 : OAI22_X1 port map( A1 => n719, A2 => n10119, B1 => n527, B2 => 
                           n10115, ZN => n7944);
   U9633 : OAI22_X1 port map( A1 => n720, A2 => n10119, B1 => n528, B2 => 
                           n10115, ZN => n7927);
   U9634 : OAI22_X1 port map( A1 => n721, A2 => n10119, B1 => n529, B2 => 
                           n10115, ZN => n7910);
   U9635 : OAI22_X1 port map( A1 => n722, A2 => n10119, B1 => n530, B2 => 
                           n10115, ZN => n7893);
   U9636 : OAI22_X1 port map( A1 => n723, A2 => n10119, B1 => n531, B2 => 
                           n10115, ZN => n7876);
   U9637 : OAI22_X1 port map( A1 => n724, A2 => n10119, B1 => n532, B2 => 
                           n10115, ZN => n7859);
   U9638 : OAI22_X1 port map( A1 => n725, A2 => n10119, B1 => n533, B2 => 
                           n10115, ZN => n7842);
   U9639 : OAI22_X1 port map( A1 => n726, A2 => n10119, B1 => n534, B2 => 
                           n10115, ZN => n7825);
   U9640 : OAI22_X1 port map( A1 => n727, A2 => n10119, B1 => n535, B2 => 
                           n10115, ZN => n7808);
   U9641 : OAI22_X1 port map( A1 => n728, A2 => n10120, B1 => n536, B2 => 
                           n10116, ZN => n7791);
   U9642 : OAI22_X1 port map( A1 => n729, A2 => n10120, B1 => n537, B2 => 
                           n10116, ZN => n7774);
   U9643 : OAI22_X1 port map( A1 => n730, A2 => n10120, B1 => n538, B2 => 
                           n10116, ZN => n7757);
   U9644 : OAI22_X1 port map( A1 => n731, A2 => n10120, B1 => n539, B2 => 
                           n10116, ZN => n7740);
   U9645 : OAI22_X1 port map( A1 => n732, A2 => n10120, B1 => n540, B2 => 
                           n10116, ZN => n7723);
   U9646 : OAI22_X1 port map( A1 => n733, A2 => n10120, B1 => n541, B2 => 
                           n10116, ZN => n7706);
   U9647 : OAI22_X1 port map( A1 => n734, A2 => n10120, B1 => n542, B2 => 
                           n10116, ZN => n7689);
   U9648 : OAI22_X1 port map( A1 => n735, A2 => n10120, B1 => n543, B2 => 
                           n10116, ZN => n7640);
   U9649 : OAI22_X1 port map( A1 => n10132, A2 => n9749, B1 => n7544, B2 => 
                           n9745, ZN => n1344);
   U9650 : OAI22_X1 port map( A1 => n10135, A2 => n9749, B1 => n7543, B2 => 
                           n9745, ZN => n1345);
   U9651 : OAI22_X1 port map( A1 => n10138, A2 => n9749, B1 => n7542, B2 => 
                           n9745, ZN => n1346);
   U9652 : OAI22_X1 port map( A1 => n10141, A2 => n9749, B1 => n7541, B2 => 
                           n9745, ZN => n1347);
   U9653 : OAI22_X1 port map( A1 => n10144, A2 => n9749, B1 => n7540, B2 => 
                           n9745, ZN => n1348);
   U9654 : OAI22_X1 port map( A1 => n10147, A2 => n9749, B1 => n7539, B2 => 
                           n9745, ZN => n1349);
   U9655 : OAI22_X1 port map( A1 => n10150, A2 => n9749, B1 => n7538, B2 => 
                           n9745, ZN => n1350);
   U9656 : OAI22_X1 port map( A1 => n10153, A2 => n9749, B1 => n7537, B2 => 
                           n9745, ZN => n1351);
   U9657 : OAI22_X1 port map( A1 => n10156, A2 => n9749, B1 => n7536, B2 => 
                           n9745, ZN => n1352);
   U9658 : OAI22_X1 port map( A1 => n10159, A2 => n9749, B1 => n7535, B2 => 
                           n9745, ZN => n1353);
   U9659 : OAI22_X1 port map( A1 => n10162, A2 => n9749, B1 => n7534, B2 => 
                           n9745, ZN => n1354);
   U9660 : OAI22_X1 port map( A1 => n10165, A2 => n9750, B1 => n7533, B2 => 
                           n9745, ZN => n1355);
   U9661 : OAI22_X1 port map( A1 => n10168, A2 => n9750, B1 => n7532, B2 => 
                           n9746, ZN => n1356);
   U9662 : OAI22_X1 port map( A1 => n10171, A2 => n9750, B1 => n7531, B2 => 
                           n9746, ZN => n1357);
   U9663 : OAI22_X1 port map( A1 => n10174, A2 => n9750, B1 => n7530, B2 => 
                           n9746, ZN => n1358);
   U9664 : OAI22_X1 port map( A1 => n10177, A2 => n9750, B1 => n7529, B2 => 
                           n9746, ZN => n1359);
   U9665 : OAI22_X1 port map( A1 => n10180, A2 => n9750, B1 => n7528, B2 => 
                           n9746, ZN => n1360);
   U9666 : OAI22_X1 port map( A1 => n10183, A2 => n9750, B1 => n7527, B2 => 
                           n9746, ZN => n1361);
   U9667 : OAI22_X1 port map( A1 => n10186, A2 => n9750, B1 => n7526, B2 => 
                           n9746, ZN => n1362);
   U9668 : OAI22_X1 port map( A1 => n10189, A2 => n9750, B1 => n7525, B2 => 
                           n9746, ZN => n1363);
   U9669 : OAI22_X1 port map( A1 => n10192, A2 => n9750, B1 => n7524, B2 => 
                           n9746, ZN => n1364);
   U9670 : OAI22_X1 port map( A1 => n10195, A2 => n9750, B1 => n7523, B2 => 
                           n9746, ZN => n1365);
   U9671 : OAI22_X1 port map( A1 => n10198, A2 => n9750, B1 => n7522, B2 => 
                           n9746, ZN => n1366);
   U9672 : OAI22_X1 port map( A1 => n10201, A2 => n9751, B1 => n7521, B2 => 
                           n9746, ZN => n1367);
   U9673 : OAI22_X1 port map( A1 => n10204, A2 => n9751, B1 => n7496, B2 => 
                           n9747, ZN => n1368);
   U9674 : OAI22_X1 port map( A1 => n10207, A2 => n9751, B1 => n7495, B2 => 
                           n9747, ZN => n1369);
   U9675 : OAI22_X1 port map( A1 => n10210, A2 => n9751, B1 => n7494, B2 => 
                           n9747, ZN => n1370);
   U9676 : OAI22_X1 port map( A1 => n10213, A2 => n9751, B1 => n7493, B2 => 
                           n9747, ZN => n1371);
   U9677 : OAI22_X1 port map( A1 => n10216, A2 => n9751, B1 => n7492, B2 => 
                           n9747, ZN => n1372);
   U9678 : OAI22_X1 port map( A1 => n10219, A2 => n9751, B1 => n7491, B2 => 
                           n9747, ZN => n1373);
   U9679 : OAI22_X1 port map( A1 => n10222, A2 => n9751, B1 => n7490, B2 => 
                           n9747, ZN => n1374);
   U9680 : OAI22_X1 port map( A1 => n10225, A2 => n9751, B1 => n7489, B2 => 
                           n9747, ZN => n1375);
   U9681 : OAI22_X1 port map( A1 => n10132, A2 => n9741, B1 => n7488, B2 => 
                           n9737, ZN => n1312);
   U9682 : OAI22_X1 port map( A1 => n10135, A2 => n9741, B1 => n7487, B2 => 
                           n9737, ZN => n1313);
   U9683 : OAI22_X1 port map( A1 => n10138, A2 => n9741, B1 => n7486, B2 => 
                           n9737, ZN => n1314);
   U9684 : OAI22_X1 port map( A1 => n10141, A2 => n9741, B1 => n7485, B2 => 
                           n9737, ZN => n1315);
   U9685 : OAI22_X1 port map( A1 => n10144, A2 => n9741, B1 => n7484, B2 => 
                           n9737, ZN => n1316);
   U9686 : OAI22_X1 port map( A1 => n10147, A2 => n9741, B1 => n7483, B2 => 
                           n9737, ZN => n1317);
   U9687 : OAI22_X1 port map( A1 => n10150, A2 => n9741, B1 => n7482, B2 => 
                           n9737, ZN => n1318);
   U9688 : OAI22_X1 port map( A1 => n10153, A2 => n9741, B1 => n7481, B2 => 
                           n9737, ZN => n1319);
   U9689 : OAI22_X1 port map( A1 => n10156, A2 => n9741, B1 => n7480, B2 => 
                           n9737, ZN => n1320);
   U9690 : OAI22_X1 port map( A1 => n10159, A2 => n9741, B1 => n7479, B2 => 
                           n9737, ZN => n1321);
   U9691 : OAI22_X1 port map( A1 => n10162, A2 => n9741, B1 => n7478, B2 => 
                           n9737, ZN => n1322);
   U9692 : OAI22_X1 port map( A1 => n10165, A2 => n9742, B1 => n7477, B2 => 
                           n9737, ZN => n1323);
   U9693 : OAI22_X1 port map( A1 => n10168, A2 => n9742, B1 => n7476, B2 => 
                           n9738, ZN => n1324);
   U9694 : OAI22_X1 port map( A1 => n10171, A2 => n9742, B1 => n7475, B2 => 
                           n9738, ZN => n1325);
   U9695 : OAI22_X1 port map( A1 => n10174, A2 => n9742, B1 => n7474, B2 => 
                           n9738, ZN => n1326);
   U9696 : OAI22_X1 port map( A1 => n10177, A2 => n9742, B1 => n7473, B2 => 
                           n9738, ZN => n1327);
   U9697 : OAI22_X1 port map( A1 => n10180, A2 => n9742, B1 => n7472, B2 => 
                           n9738, ZN => n1328);
   U9698 : OAI22_X1 port map( A1 => n10183, A2 => n9742, B1 => n7471, B2 => 
                           n9738, ZN => n1329);
   U9699 : OAI22_X1 port map( A1 => n10186, A2 => n9742, B1 => n7470, B2 => 
                           n9738, ZN => n1330);
   U9700 : OAI22_X1 port map( A1 => n10189, A2 => n9742, B1 => n7469, B2 => 
                           n9738, ZN => n1331);
   U9701 : OAI22_X1 port map( A1 => n10192, A2 => n9742, B1 => n7468, B2 => 
                           n9738, ZN => n1332);
   U9702 : OAI22_X1 port map( A1 => n10195, A2 => n9742, B1 => n7467, B2 => 
                           n9738, ZN => n1333);
   U9703 : OAI22_X1 port map( A1 => n10198, A2 => n9742, B1 => n7466, B2 => 
                           n9738, ZN => n1334);
   U9704 : OAI22_X1 port map( A1 => n10201, A2 => n9743, B1 => n7465, B2 => 
                           n9738, ZN => n1335);
   U9705 : OAI22_X1 port map( A1 => n10204, A2 => n9743, B1 => n7464, B2 => 
                           n9739, ZN => n1336);
   U9706 : OAI22_X1 port map( A1 => n10207, A2 => n9743, B1 => n7463, B2 => 
                           n9739, ZN => n1337);
   U9707 : OAI22_X1 port map( A1 => n10210, A2 => n9743, B1 => n7462, B2 => 
                           n9739, ZN => n1338);
   U9708 : OAI22_X1 port map( A1 => n10213, A2 => n9743, B1 => n7461, B2 => 
                           n9739, ZN => n1339);
   U9709 : OAI22_X1 port map( A1 => n10216, A2 => n9743, B1 => n7460, B2 => 
                           n9739, ZN => n1340);
   U9710 : OAI22_X1 port map( A1 => n10219, A2 => n9743, B1 => n7459, B2 => 
                           n9739, ZN => n1341);
   U9711 : OAI22_X1 port map( A1 => n10222, A2 => n9743, B1 => n7458, B2 => 
                           n9739, ZN => n1342);
   U9712 : OAI22_X1 port map( A1 => n10225, A2 => n9743, B1 => n7457, B2 => 
                           n9739, ZN => n1343);
   U9713 : OAI22_X1 port map( A1 => n10131, A2 => n9853, B1 => n7328, B2 => 
                           n9849, ZN => n1760);
   U9714 : OAI22_X1 port map( A1 => n10134, A2 => n9853, B1 => n7327, B2 => 
                           n9849, ZN => n1761);
   U9715 : OAI22_X1 port map( A1 => n10137, A2 => n9853, B1 => n7326, B2 => 
                           n9849, ZN => n1762);
   U9716 : OAI22_X1 port map( A1 => n10140, A2 => n9853, B1 => n7325, B2 => 
                           n9849, ZN => n1763);
   U9717 : OAI22_X1 port map( A1 => n10143, A2 => n9853, B1 => n7324, B2 => 
                           n9849, ZN => n1764);
   U9718 : OAI22_X1 port map( A1 => n10146, A2 => n9853, B1 => n7323, B2 => 
                           n9849, ZN => n1765);
   U9719 : OAI22_X1 port map( A1 => n10149, A2 => n9853, B1 => n7322, B2 => 
                           n9849, ZN => n1766);
   U9720 : OAI22_X1 port map( A1 => n10152, A2 => n9853, B1 => n7321, B2 => 
                           n9849, ZN => n1767);
   U9721 : OAI22_X1 port map( A1 => n10155, A2 => n9853, B1 => n7320, B2 => 
                           n9849, ZN => n1768);
   U9722 : OAI22_X1 port map( A1 => n10158, A2 => n9853, B1 => n7319, B2 => 
                           n9849, ZN => n1769);
   U9723 : OAI22_X1 port map( A1 => n10161, A2 => n9853, B1 => n7318, B2 => 
                           n9849, ZN => n1770);
   U9724 : OAI22_X1 port map( A1 => n10164, A2 => n9854, B1 => n7317, B2 => 
                           n9849, ZN => n1771);
   U9725 : OAI22_X1 port map( A1 => n10167, A2 => n9854, B1 => n7316, B2 => 
                           n9850, ZN => n1772);
   U9726 : OAI22_X1 port map( A1 => n10170, A2 => n9854, B1 => n7315, B2 => 
                           n9850, ZN => n1773);
   U9727 : OAI22_X1 port map( A1 => n10173, A2 => n9854, B1 => n7314, B2 => 
                           n9850, ZN => n1774);
   U9728 : OAI22_X1 port map( A1 => n10176, A2 => n9854, B1 => n7313, B2 => 
                           n9850, ZN => n1775);
   U9729 : OAI22_X1 port map( A1 => n10179, A2 => n9854, B1 => n7312, B2 => 
                           n9850, ZN => n1776);
   U9730 : OAI22_X1 port map( A1 => n10182, A2 => n9854, B1 => n7311, B2 => 
                           n9850, ZN => n1777);
   U9731 : OAI22_X1 port map( A1 => n10185, A2 => n9854, B1 => n7310, B2 => 
                           n9850, ZN => n1778);
   U9732 : OAI22_X1 port map( A1 => n10188, A2 => n9854, B1 => n7309, B2 => 
                           n9850, ZN => n1779);
   U9733 : OAI22_X1 port map( A1 => n10191, A2 => n9854, B1 => n7308, B2 => 
                           n9850, ZN => n1780);
   U9734 : OAI22_X1 port map( A1 => n10194, A2 => n9854, B1 => n7307, B2 => 
                           n9850, ZN => n1781);
   U9735 : OAI22_X1 port map( A1 => n10197, A2 => n9854, B1 => n7306, B2 => 
                           n9850, ZN => n1782);
   U9736 : OAI22_X1 port map( A1 => n10200, A2 => n9855, B1 => n7305, B2 => 
                           n9850, ZN => n1783);
   U9737 : OAI22_X1 port map( A1 => n10203, A2 => n9855, B1 => n7304, B2 => 
                           n9851, ZN => n1784);
   U9738 : OAI22_X1 port map( A1 => n10206, A2 => n9855, B1 => n7303, B2 => 
                           n9851, ZN => n1785);
   U9739 : OAI22_X1 port map( A1 => n10209, A2 => n9855, B1 => n7302, B2 => 
                           n9851, ZN => n1786);
   U9740 : OAI22_X1 port map( A1 => n10212, A2 => n9855, B1 => n7301, B2 => 
                           n9851, ZN => n1787);
   U9741 : OAI22_X1 port map( A1 => n10215, A2 => n9855, B1 => n7300, B2 => 
                           n9851, ZN => n1788);
   U9742 : OAI22_X1 port map( A1 => n10218, A2 => n9855, B1 => n7299, B2 => 
                           n9851, ZN => n1789);
   U9743 : OAI22_X1 port map( A1 => n10221, A2 => n9855, B1 => n7298, B2 => 
                           n9851, ZN => n1790);
   U9744 : OAI22_X1 port map( A1 => n10224, A2 => n9855, B1 => n7297, B2 => 
                           n9851, ZN => n1791);
   U9745 : OAI22_X1 port map( A1 => n10130, A2 => n9893, B1 => n7201, B2 => 
                           n9889, ZN => n1920);
   U9746 : OAI22_X1 port map( A1 => n10133, A2 => n9893, B1 => n7200, B2 => 
                           n9889, ZN => n1921);
   U9747 : OAI22_X1 port map( A1 => n10136, A2 => n9893, B1 => n7199, B2 => 
                           n9889, ZN => n1922);
   U9748 : OAI22_X1 port map( A1 => n10139, A2 => n9893, B1 => n7198, B2 => 
                           n9889, ZN => n1923);
   U9749 : OAI22_X1 port map( A1 => n10142, A2 => n9893, B1 => n7197, B2 => 
                           n9889, ZN => n1924);
   U9750 : OAI22_X1 port map( A1 => n10145, A2 => n9893, B1 => n7196, B2 => 
                           n9889, ZN => n1925);
   U9751 : OAI22_X1 port map( A1 => n10148, A2 => n9893, B1 => n7195, B2 => 
                           n9889, ZN => n1926);
   U9752 : OAI22_X1 port map( A1 => n10151, A2 => n9893, B1 => n7194, B2 => 
                           n9889, ZN => n1927);
   U9753 : OAI22_X1 port map( A1 => n10154, A2 => n9893, B1 => n7193, B2 => 
                           n9889, ZN => n1928);
   U9754 : OAI22_X1 port map( A1 => n10157, A2 => n9893, B1 => n7192, B2 => 
                           n9889, ZN => n1929);
   U9755 : OAI22_X1 port map( A1 => n10160, A2 => n9893, B1 => n7191, B2 => 
                           n9889, ZN => n1930);
   U9756 : OAI22_X1 port map( A1 => n10163, A2 => n9894, B1 => n7190, B2 => 
                           n9889, ZN => n1931);
   U9757 : OAI22_X1 port map( A1 => n10166, A2 => n9894, B1 => n7189, B2 => 
                           n9890, ZN => n1932);
   U9758 : OAI22_X1 port map( A1 => n10169, A2 => n9894, B1 => n7188, B2 => 
                           n9890, ZN => n1933);
   U9759 : OAI22_X1 port map( A1 => n10172, A2 => n9894, B1 => n7187, B2 => 
                           n9890, ZN => n1934);
   U9760 : OAI22_X1 port map( A1 => n10175, A2 => n9894, B1 => n7186, B2 => 
                           n9890, ZN => n1935);
   U9761 : OAI22_X1 port map( A1 => n10178, A2 => n9894, B1 => n7185, B2 => 
                           n9890, ZN => n1936);
   U9762 : OAI22_X1 port map( A1 => n10181, A2 => n9894, B1 => n7184, B2 => 
                           n9890, ZN => n1937);
   U9763 : OAI22_X1 port map( A1 => n10184, A2 => n9894, B1 => n7183, B2 => 
                           n9890, ZN => n1938);
   U9764 : OAI22_X1 port map( A1 => n10187, A2 => n9894, B1 => n7182, B2 => 
                           n9890, ZN => n1939);
   U9765 : OAI22_X1 port map( A1 => n10190, A2 => n9894, B1 => n7181, B2 => 
                           n9890, ZN => n1940);
   U9766 : OAI22_X1 port map( A1 => n10193, A2 => n9894, B1 => n7180, B2 => 
                           n9890, ZN => n1941);
   U9767 : OAI22_X1 port map( A1 => n10196, A2 => n9894, B1 => n7179, B2 => 
                           n9890, ZN => n1942);
   U9768 : OAI22_X1 port map( A1 => n10199, A2 => n9895, B1 => n7178, B2 => 
                           n9890, ZN => n1943);
   U9769 : OAI22_X1 port map( A1 => n10202, A2 => n9895, B1 => n7177, B2 => 
                           n9891, ZN => n1944);
   U9770 : OAI22_X1 port map( A1 => n10205, A2 => n9895, B1 => n7176, B2 => 
                           n9891, ZN => n1945);
   U9771 : OAI22_X1 port map( A1 => n10208, A2 => n9895, B1 => n7175, B2 => 
                           n9891, ZN => n1946);
   U9772 : OAI22_X1 port map( A1 => n10211, A2 => n9895, B1 => n7174, B2 => 
                           n9891, ZN => n1947);
   U9773 : OAI22_X1 port map( A1 => n10214, A2 => n9895, B1 => n7173, B2 => 
                           n9891, ZN => n1948);
   U9774 : OAI22_X1 port map( A1 => n10217, A2 => n9895, B1 => n7172, B2 => 
                           n9891, ZN => n1949);
   U9775 : OAI22_X1 port map( A1 => n10220, A2 => n9895, B1 => n7171, B2 => 
                           n9891, ZN => n1950);
   U9776 : OAI22_X1 port map( A1 => n10223, A2 => n9895, B1 => n7170, B2 => 
                           n9891, ZN => n1951);
   U9777 : OAI22_X1 port map( A1 => n10130, A2 => n9901, B1 => n7169, B2 => 
                           n9897, ZN => n1952);
   U9778 : OAI22_X1 port map( A1 => n10133, A2 => n9901, B1 => n7168, B2 => 
                           n9897, ZN => n1953);
   U9779 : OAI22_X1 port map( A1 => n10136, A2 => n9901, B1 => n7167, B2 => 
                           n9897, ZN => n1954);
   U9780 : OAI22_X1 port map( A1 => n10139, A2 => n9901, B1 => n7166, B2 => 
                           n9897, ZN => n1955);
   U9781 : OAI22_X1 port map( A1 => n10142, A2 => n9901, B1 => n7165, B2 => 
                           n9897, ZN => n1956);
   U9782 : OAI22_X1 port map( A1 => n10145, A2 => n9901, B1 => n7164, B2 => 
                           n9897, ZN => n1957);
   U9783 : OAI22_X1 port map( A1 => n10148, A2 => n9901, B1 => n7163, B2 => 
                           n9897, ZN => n1958);
   U9784 : OAI22_X1 port map( A1 => n10151, A2 => n9901, B1 => n7162, B2 => 
                           n9897, ZN => n1959);
   U9785 : OAI22_X1 port map( A1 => n10154, A2 => n9901, B1 => n7161, B2 => 
                           n9897, ZN => n1960);
   U9786 : OAI22_X1 port map( A1 => n10157, A2 => n9901, B1 => n7160, B2 => 
                           n9897, ZN => n1961);
   U9787 : OAI22_X1 port map( A1 => n10160, A2 => n9901, B1 => n7159, B2 => 
                           n9897, ZN => n1962);
   U9788 : OAI22_X1 port map( A1 => n10163, A2 => n9902, B1 => n7158, B2 => 
                           n9897, ZN => n1963);
   U9789 : OAI22_X1 port map( A1 => n10166, A2 => n9902, B1 => n7157, B2 => 
                           n9898, ZN => n1964);
   U9790 : OAI22_X1 port map( A1 => n10169, A2 => n9902, B1 => n7156, B2 => 
                           n9898, ZN => n1965);
   U9791 : OAI22_X1 port map( A1 => n10172, A2 => n9902, B1 => n7155, B2 => 
                           n9898, ZN => n1966);
   U9792 : OAI22_X1 port map( A1 => n10175, A2 => n9902, B1 => n7154, B2 => 
                           n9898, ZN => n1967);
   U9793 : OAI22_X1 port map( A1 => n10178, A2 => n9902, B1 => n7153, B2 => 
                           n9898, ZN => n1968);
   U9794 : OAI22_X1 port map( A1 => n10181, A2 => n9902, B1 => n7152, B2 => 
                           n9898, ZN => n1969);
   U9795 : OAI22_X1 port map( A1 => n10184, A2 => n9902, B1 => n7151, B2 => 
                           n9898, ZN => n1970);
   U9796 : OAI22_X1 port map( A1 => n10187, A2 => n9902, B1 => n7150, B2 => 
                           n9898, ZN => n1971);
   U9797 : OAI22_X1 port map( A1 => n10190, A2 => n9902, B1 => n7149, B2 => 
                           n9898, ZN => n1972);
   U9798 : OAI22_X1 port map( A1 => n10193, A2 => n9902, B1 => n7148, B2 => 
                           n9898, ZN => n1973);
   U9799 : OAI22_X1 port map( A1 => n10196, A2 => n9902, B1 => n7147, B2 => 
                           n9898, ZN => n1974);
   U9800 : OAI22_X1 port map( A1 => n10199, A2 => n9903, B1 => n7146, B2 => 
                           n9898, ZN => n1975);
   U9801 : OAI22_X1 port map( A1 => n10202, A2 => n9903, B1 => n7145, B2 => 
                           n9899, ZN => n1976);
   U9802 : OAI22_X1 port map( A1 => n10205, A2 => n9903, B1 => n7144, B2 => 
                           n9899, ZN => n1977);
   U9803 : OAI22_X1 port map( A1 => n10208, A2 => n9903, B1 => n7143, B2 => 
                           n9899, ZN => n1978);
   U9804 : OAI22_X1 port map( A1 => n10211, A2 => n9903, B1 => n7142, B2 => 
                           n9899, ZN => n1979);
   U9805 : OAI22_X1 port map( A1 => n10214, A2 => n9903, B1 => n7141, B2 => 
                           n9899, ZN => n1980);
   U9806 : OAI22_X1 port map( A1 => n10217, A2 => n9903, B1 => n7140, B2 => 
                           n9899, ZN => n1981);
   U9807 : OAI22_X1 port map( A1 => n10220, A2 => n9903, B1 => n7139, B2 => 
                           n9899, ZN => n1982);
   U9808 : OAI22_X1 port map( A1 => n10223, A2 => n9903, B1 => n7138, B2 => 
                           n9899, ZN => n1983);
   U9809 : OAI22_X1 port map( A1 => n10130, A2 => n9973, B1 => n6881, B2 => 
                           n9969, ZN => n2240);
   U9810 : OAI22_X1 port map( A1 => n10133, A2 => n9973, B1 => n6880, B2 => 
                           n9969, ZN => n2241);
   U9811 : OAI22_X1 port map( A1 => n10136, A2 => n9973, B1 => n6879, B2 => 
                           n9969, ZN => n2242);
   U9812 : OAI22_X1 port map( A1 => n10139, A2 => n9973, B1 => n6878, B2 => 
                           n9969, ZN => n2243);
   U9813 : OAI22_X1 port map( A1 => n10142, A2 => n9973, B1 => n6877, B2 => 
                           n9969, ZN => n2244);
   U9814 : OAI22_X1 port map( A1 => n10145, A2 => n9973, B1 => n6876, B2 => 
                           n9969, ZN => n2245);
   U9815 : OAI22_X1 port map( A1 => n10148, A2 => n9973, B1 => n6875, B2 => 
                           n9969, ZN => n2246);
   U9816 : OAI22_X1 port map( A1 => n10151, A2 => n9973, B1 => n6874, B2 => 
                           n9969, ZN => n2247);
   U9817 : OAI22_X1 port map( A1 => n10154, A2 => n9973, B1 => n6873, B2 => 
                           n9969, ZN => n2248);
   U9818 : OAI22_X1 port map( A1 => n10157, A2 => n9973, B1 => n6872, B2 => 
                           n9969, ZN => n2249);
   U9819 : OAI22_X1 port map( A1 => n10160, A2 => n9973, B1 => n6871, B2 => 
                           n9969, ZN => n2250);
   U9820 : OAI22_X1 port map( A1 => n10163, A2 => n9974, B1 => n6870, B2 => 
                           n9969, ZN => n2251);
   U9821 : OAI22_X1 port map( A1 => n10166, A2 => n9974, B1 => n6869, B2 => 
                           n9970, ZN => n2252);
   U9822 : OAI22_X1 port map( A1 => n10169, A2 => n9974, B1 => n6868, B2 => 
                           n9970, ZN => n2253);
   U9823 : OAI22_X1 port map( A1 => n10172, A2 => n9974, B1 => n6867, B2 => 
                           n9970, ZN => n2254);
   U9824 : OAI22_X1 port map( A1 => n10175, A2 => n9974, B1 => n6866, B2 => 
                           n9970, ZN => n2255);
   U9825 : OAI22_X1 port map( A1 => n10178, A2 => n9974, B1 => n6865, B2 => 
                           n9970, ZN => n2256);
   U9826 : OAI22_X1 port map( A1 => n10181, A2 => n9974, B1 => n6864, B2 => 
                           n9970, ZN => n2257);
   U9827 : OAI22_X1 port map( A1 => n10184, A2 => n9974, B1 => n6863, B2 => 
                           n9970, ZN => n2258);
   U9828 : OAI22_X1 port map( A1 => n10187, A2 => n9974, B1 => n6862, B2 => 
                           n9970, ZN => n2259);
   U9829 : OAI22_X1 port map( A1 => n10190, A2 => n9974, B1 => n6861, B2 => 
                           n9970, ZN => n2260);
   U9830 : OAI22_X1 port map( A1 => n10193, A2 => n9974, B1 => n6860, B2 => 
                           n9970, ZN => n2261);
   U9831 : OAI22_X1 port map( A1 => n10196, A2 => n9974, B1 => n6859, B2 => 
                           n9970, ZN => n2262);
   U9832 : OAI22_X1 port map( A1 => n10199, A2 => n9975, B1 => n6858, B2 => 
                           n9970, ZN => n2263);
   U9833 : OAI22_X1 port map( A1 => n10202, A2 => n9975, B1 => n6857, B2 => 
                           n9971, ZN => n2264);
   U9834 : OAI22_X1 port map( A1 => n10205, A2 => n9975, B1 => n6856, B2 => 
                           n9971, ZN => n2265);
   U9835 : OAI22_X1 port map( A1 => n10208, A2 => n9975, B1 => n6855, B2 => 
                           n9971, ZN => n2266);
   U9836 : OAI22_X1 port map( A1 => n10211, A2 => n9975, B1 => n6854, B2 => 
                           n9971, ZN => n2267);
   U9837 : OAI22_X1 port map( A1 => n10214, A2 => n9975, B1 => n6853, B2 => 
                           n9971, ZN => n2268);
   U9838 : OAI22_X1 port map( A1 => n10217, A2 => n9975, B1 => n6852, B2 => 
                           n9971, ZN => n2269);
   U9839 : OAI22_X1 port map( A1 => n10220, A2 => n9975, B1 => n6851, B2 => 
                           n9971, ZN => n2270);
   U9840 : OAI22_X1 port map( A1 => n10223, A2 => n9975, B1 => n6850, B2 => 
                           n9971, ZN => n2271);
   U9841 : OAI22_X1 port map( A1 => n10130, A2 => n9981, B1 => n6849, B2 => 
                           n9977, ZN => n2272);
   U9842 : OAI22_X1 port map( A1 => n10133, A2 => n9981, B1 => n6848, B2 => 
                           n9977, ZN => n2273);
   U9843 : OAI22_X1 port map( A1 => n10136, A2 => n9981, B1 => n6847, B2 => 
                           n9977, ZN => n2274);
   U9844 : OAI22_X1 port map( A1 => n10139, A2 => n9981, B1 => n6846, B2 => 
                           n9977, ZN => n2275);
   U9845 : OAI22_X1 port map( A1 => n10142, A2 => n9981, B1 => n6845, B2 => 
                           n9977, ZN => n2276);
   U9846 : OAI22_X1 port map( A1 => n10145, A2 => n9981, B1 => n6844, B2 => 
                           n9977, ZN => n2277);
   U9847 : OAI22_X1 port map( A1 => n10148, A2 => n9981, B1 => n6843, B2 => 
                           n9977, ZN => n2278);
   U9848 : OAI22_X1 port map( A1 => n10151, A2 => n9981, B1 => n6842, B2 => 
                           n9977, ZN => n2279);
   U9849 : OAI22_X1 port map( A1 => n10154, A2 => n9981, B1 => n6841, B2 => 
                           n9977, ZN => n2280);
   U9850 : OAI22_X1 port map( A1 => n10157, A2 => n9981, B1 => n6840, B2 => 
                           n9977, ZN => n2281);
   U9851 : OAI22_X1 port map( A1 => n10160, A2 => n9981, B1 => n6839, B2 => 
                           n9977, ZN => n2282);
   U9852 : OAI22_X1 port map( A1 => n10163, A2 => n9982, B1 => n6838, B2 => 
                           n9977, ZN => n2283);
   U9853 : OAI22_X1 port map( A1 => n10166, A2 => n9982, B1 => n6837, B2 => 
                           n9978, ZN => n2284);
   U9854 : OAI22_X1 port map( A1 => n10169, A2 => n9982, B1 => n6836, B2 => 
                           n9978, ZN => n2285);
   U9855 : OAI22_X1 port map( A1 => n10172, A2 => n9982, B1 => n6835, B2 => 
                           n9978, ZN => n2286);
   U9856 : OAI22_X1 port map( A1 => n10175, A2 => n9982, B1 => n6834, B2 => 
                           n9978, ZN => n2287);
   U9857 : OAI22_X1 port map( A1 => n10178, A2 => n9982, B1 => n6833, B2 => 
                           n9978, ZN => n2288);
   U9858 : OAI22_X1 port map( A1 => n10181, A2 => n9982, B1 => n6832, B2 => 
                           n9978, ZN => n2289);
   U9859 : OAI22_X1 port map( A1 => n10184, A2 => n9982, B1 => n6831, B2 => 
                           n9978, ZN => n2290);
   U9860 : OAI22_X1 port map( A1 => n10187, A2 => n9982, B1 => n6830, B2 => 
                           n9978, ZN => n2291);
   U9861 : OAI22_X1 port map( A1 => n10190, A2 => n9982, B1 => n6829, B2 => 
                           n9978, ZN => n2292);
   U9862 : OAI22_X1 port map( A1 => n10193, A2 => n9982, B1 => n6828, B2 => 
                           n9978, ZN => n2293);
   U9863 : OAI22_X1 port map( A1 => n10196, A2 => n9982, B1 => n6827, B2 => 
                           n9978, ZN => n2294);
   U9864 : OAI22_X1 port map( A1 => n10199, A2 => n9983, B1 => n6826, B2 => 
                           n9978, ZN => n2295);
   U9865 : OAI22_X1 port map( A1 => n10202, A2 => n9983, B1 => n6825, B2 => 
                           n9979, ZN => n2296);
   U9866 : OAI22_X1 port map( A1 => n10205, A2 => n9983, B1 => n6824, B2 => 
                           n9979, ZN => n2297);
   U9867 : OAI22_X1 port map( A1 => n10208, A2 => n9983, B1 => n6823, B2 => 
                           n9979, ZN => n2298);
   U9868 : OAI22_X1 port map( A1 => n10211, A2 => n9983, B1 => n6822, B2 => 
                           n9979, ZN => n2299);
   U9869 : OAI22_X1 port map( A1 => n10214, A2 => n9983, B1 => n6821, B2 => 
                           n9979, ZN => n2300);
   U9870 : OAI22_X1 port map( A1 => n10217, A2 => n9983, B1 => n6820, B2 => 
                           n9979, ZN => n2301);
   U9871 : OAI22_X1 port map( A1 => n10220, A2 => n9983, B1 => n6819, B2 => 
                           n9979, ZN => n2302);
   U9872 : OAI22_X1 port map( A1 => n10223, A2 => n9983, B1 => n6818, B2 => 
                           n9979, ZN => n2303);
   U9873 : OAI22_X1 port map( A1 => n10224, A2 => n9871, B1 => n7633, B2 => 
                           n9867, ZN => n1855);
   U9874 : OAI22_X1 port map( A1 => n10132, A2 => n9781, B1 => n7592, B2 => 
                           n9777, ZN => n1472);
   U9875 : OAI22_X1 port map( A1 => n10135, A2 => n9781, B1 => n7591, B2 => 
                           n9777, ZN => n1473);
   U9876 : OAI22_X1 port map( A1 => n10138, A2 => n9781, B1 => n7590, B2 => 
                           n9777, ZN => n1474);
   U9877 : OAI22_X1 port map( A1 => n10141, A2 => n9781, B1 => n7589, B2 => 
                           n9777, ZN => n1475);
   U9878 : OAI22_X1 port map( A1 => n10144, A2 => n9781, B1 => n7588, B2 => 
                           n9777, ZN => n1476);
   U9879 : OAI22_X1 port map( A1 => n10147, A2 => n9781, B1 => n7587, B2 => 
                           n9777, ZN => n1477);
   U9880 : OAI22_X1 port map( A1 => n10150, A2 => n9781, B1 => n7586, B2 => 
                           n9777, ZN => n1478);
   U9881 : OAI22_X1 port map( A1 => n10153, A2 => n9781, B1 => n7585, B2 => 
                           n9777, ZN => n1479);
   U9882 : OAI22_X1 port map( A1 => n10156, A2 => n9781, B1 => n7584, B2 => 
                           n9777, ZN => n1480);
   U9883 : OAI22_X1 port map( A1 => n10159, A2 => n9781, B1 => n7583, B2 => 
                           n9777, ZN => n1481);
   U9884 : OAI22_X1 port map( A1 => n10162, A2 => n9781, B1 => n7582, B2 => 
                           n9777, ZN => n1482);
   U9885 : OAI22_X1 port map( A1 => n10165, A2 => n9782, B1 => n7581, B2 => 
                           n9777, ZN => n1483);
   U9886 : OAI22_X1 port map( A1 => n10168, A2 => n9782, B1 => n7580, B2 => 
                           n9778, ZN => n1484);
   U9887 : OAI22_X1 port map( A1 => n10171, A2 => n9782, B1 => n7579, B2 => 
                           n9778, ZN => n1485);
   U9888 : OAI22_X1 port map( A1 => n10174, A2 => n9782, B1 => n7578, B2 => 
                           n9778, ZN => n1486);
   U9889 : OAI22_X1 port map( A1 => n10177, A2 => n9782, B1 => n7577, B2 => 
                           n9778, ZN => n1487);
   U9890 : OAI22_X1 port map( A1 => n10180, A2 => n9782, B1 => n7576, B2 => 
                           n9778, ZN => n1488);
   U9891 : OAI22_X1 port map( A1 => n10183, A2 => n9782, B1 => n7575, B2 => 
                           n9778, ZN => n1489);
   U9892 : OAI22_X1 port map( A1 => n10186, A2 => n9782, B1 => n7574, B2 => 
                           n9778, ZN => n1490);
   U9893 : OAI22_X1 port map( A1 => n10189, A2 => n9782, B1 => n7573, B2 => 
                           n9778, ZN => n1491);
   U9894 : OAI22_X1 port map( A1 => n10192, A2 => n9782, B1 => n7572, B2 => 
                           n9778, ZN => n1492);
   U9895 : OAI22_X1 port map( A1 => n10195, A2 => n9782, B1 => n7571, B2 => 
                           n9778, ZN => n1493);
   U9896 : OAI22_X1 port map( A1 => n10198, A2 => n9782, B1 => n7570, B2 => 
                           n9778, ZN => n1494);
   U9897 : OAI22_X1 port map( A1 => n10201, A2 => n9783, B1 => n7569, B2 => 
                           n9778, ZN => n1495);
   U9898 : OAI22_X1 port map( A1 => n10132, A2 => n9757, B1 => n7568, B2 => 
                           n9753, ZN => n1376);
   U9899 : OAI22_X1 port map( A1 => n10135, A2 => n9757, B1 => n7567, B2 => 
                           n9753, ZN => n1377);
   U9900 : OAI22_X1 port map( A1 => n10138, A2 => n9757, B1 => n7566, B2 => 
                           n9753, ZN => n1378);
   U9901 : OAI22_X1 port map( A1 => n10141, A2 => n9757, B1 => n7565, B2 => 
                           n9753, ZN => n1379);
   U9902 : OAI22_X1 port map( A1 => n10144, A2 => n9757, B1 => n7564, B2 => 
                           n9753, ZN => n1380);
   U9903 : OAI22_X1 port map( A1 => n10147, A2 => n9757, B1 => n7563, B2 => 
                           n9753, ZN => n1381);
   U9904 : OAI22_X1 port map( A1 => n10150, A2 => n9757, B1 => n7562, B2 => 
                           n9753, ZN => n1382);
   U9905 : OAI22_X1 port map( A1 => n10153, A2 => n9757, B1 => n7561, B2 => 
                           n9753, ZN => n1383);
   U9906 : OAI22_X1 port map( A1 => n10156, A2 => n9757, B1 => n7560, B2 => 
                           n9753, ZN => n1384);
   U9907 : OAI22_X1 port map( A1 => n10159, A2 => n9757, B1 => n7559, B2 => 
                           n9753, ZN => n1385);
   U9908 : OAI22_X1 port map( A1 => n10162, A2 => n9757, B1 => n7558, B2 => 
                           n9753, ZN => n1386);
   U9909 : OAI22_X1 port map( A1 => n10165, A2 => n9758, B1 => n7557, B2 => 
                           n9753, ZN => n1387);
   U9910 : OAI22_X1 port map( A1 => n10168, A2 => n9758, B1 => n7556, B2 => 
                           n9754, ZN => n1388);
   U9911 : OAI22_X1 port map( A1 => n10171, A2 => n9758, B1 => n7555, B2 => 
                           n9754, ZN => n1389);
   U9912 : OAI22_X1 port map( A1 => n10174, A2 => n9758, B1 => n7554, B2 => 
                           n9754, ZN => n1390);
   U9913 : OAI22_X1 port map( A1 => n10177, A2 => n9758, B1 => n7553, B2 => 
                           n9754, ZN => n1391);
   U9914 : OAI22_X1 port map( A1 => n10180, A2 => n9758, B1 => n7552, B2 => 
                           n9754, ZN => n1392);
   U9915 : OAI22_X1 port map( A1 => n10183, A2 => n9758, B1 => n7551, B2 => 
                           n9754, ZN => n1393);
   U9916 : OAI22_X1 port map( A1 => n10186, A2 => n9758, B1 => n7550, B2 => 
                           n9754, ZN => n1394);
   U9917 : OAI22_X1 port map( A1 => n10189, A2 => n9758, B1 => n7549, B2 => 
                           n9754, ZN => n1395);
   U9918 : OAI22_X1 port map( A1 => n10192, A2 => n9758, B1 => n7548, B2 => 
                           n9754, ZN => n1396);
   U9919 : OAI22_X1 port map( A1 => n10195, A2 => n9758, B1 => n7547, B2 => 
                           n9754, ZN => n1397);
   U9920 : OAI22_X1 port map( A1 => n10198, A2 => n9758, B1 => n7546, B2 => 
                           n9754, ZN => n1398);
   U9921 : OAI22_X1 port map( A1 => n10201, A2 => n9759, B1 => n7545, B2 => 
                           n9754, ZN => n1399);
   U9922 : OAI22_X1 port map( A1 => n10204, A2 => n9783, B1 => n7512, B2 => 
                           n9779, ZN => n1496);
   U9923 : OAI22_X1 port map( A1 => n10207, A2 => n9783, B1 => n7511, B2 => 
                           n9779, ZN => n1497);
   U9924 : OAI22_X1 port map( A1 => n10210, A2 => n9783, B1 => n7510, B2 => 
                           n9779, ZN => n1498);
   U9925 : OAI22_X1 port map( A1 => n10213, A2 => n9783, B1 => n7509, B2 => 
                           n9779, ZN => n1499);
   U9926 : OAI22_X1 port map( A1 => n10216, A2 => n9783, B1 => n7508, B2 => 
                           n9779, ZN => n1500);
   U9927 : OAI22_X1 port map( A1 => n10219, A2 => n9783, B1 => n7507, B2 => 
                           n9779, ZN => n1501);
   U9928 : OAI22_X1 port map( A1 => n10222, A2 => n9783, B1 => n7506, B2 => 
                           n9779, ZN => n1502);
   U9929 : OAI22_X1 port map( A1 => n10225, A2 => n9783, B1 => n7505, B2 => 
                           n9779, ZN => n1503);
   U9930 : OAI22_X1 port map( A1 => n10204, A2 => n9759, B1 => n7504, B2 => 
                           n9755, ZN => n1400);
   U9931 : OAI22_X1 port map( A1 => n10207, A2 => n9759, B1 => n7503, B2 => 
                           n9755, ZN => n1401);
   U9932 : OAI22_X1 port map( A1 => n10210, A2 => n9759, B1 => n7502, B2 => 
                           n9755, ZN => n1402);
   U9933 : OAI22_X1 port map( A1 => n10213, A2 => n9759, B1 => n7501, B2 => 
                           n9755, ZN => n1403);
   U9934 : OAI22_X1 port map( A1 => n10216, A2 => n9759, B1 => n7500, B2 => 
                           n9755, ZN => n1404);
   U9935 : OAI22_X1 port map( A1 => n10219, A2 => n9759, B1 => n7499, B2 => 
                           n9755, ZN => n1405);
   U9936 : OAI22_X1 port map( A1 => n10222, A2 => n9759, B1 => n7498, B2 => 
                           n9755, ZN => n1406);
   U9937 : OAI22_X1 port map( A1 => n10225, A2 => n9759, B1 => n7497, B2 => 
                           n9755, ZN => n1407);
   U9938 : OAI22_X1 port map( A1 => n10131, A2 => n9869, B1 => n7296, B2 => 
                           n9865, ZN => n1824);
   U9939 : OAI22_X1 port map( A1 => n10134, A2 => n9869, B1 => n7295, B2 => 
                           n9865, ZN => n1825);
   U9940 : OAI22_X1 port map( A1 => n10137, A2 => n9869, B1 => n7294, B2 => 
                           n9865, ZN => n1826);
   U9941 : OAI22_X1 port map( A1 => n10140, A2 => n9869, B1 => n7293, B2 => 
                           n9865, ZN => n1827);
   U9942 : OAI22_X1 port map( A1 => n10143, A2 => n9869, B1 => n7292, B2 => 
                           n9865, ZN => n1828);
   U9943 : OAI22_X1 port map( A1 => n10146, A2 => n9869, B1 => n7291, B2 => 
                           n9865, ZN => n1829);
   U9944 : OAI22_X1 port map( A1 => n10149, A2 => n9869, B1 => n7290, B2 => 
                           n9865, ZN => n1830);
   U9945 : OAI22_X1 port map( A1 => n10152, A2 => n9869, B1 => n7289, B2 => 
                           n9865, ZN => n1831);
   U9946 : OAI22_X1 port map( A1 => n10155, A2 => n9869, B1 => n7288, B2 => 
                           n9865, ZN => n1832);
   U9947 : OAI22_X1 port map( A1 => n10158, A2 => n9869, B1 => n7287, B2 => 
                           n9865, ZN => n1833);
   U9948 : OAI22_X1 port map( A1 => n10161, A2 => n9869, B1 => n7286, B2 => 
                           n9865, ZN => n1834);
   U9949 : OAI22_X1 port map( A1 => n10164, A2 => n9870, B1 => n7285, B2 => 
                           n9865, ZN => n1835);
   U9950 : OAI22_X1 port map( A1 => n10167, A2 => n9870, B1 => n7284, B2 => 
                           n9866, ZN => n1836);
   U9951 : OAI22_X1 port map( A1 => n10170, A2 => n9870, B1 => n7283, B2 => 
                           n9866, ZN => n1837);
   U9952 : OAI22_X1 port map( A1 => n10173, A2 => n9870, B1 => n7282, B2 => 
                           n9866, ZN => n1838);
   U9953 : OAI22_X1 port map( A1 => n10176, A2 => n9870, B1 => n7281, B2 => 
                           n9866, ZN => n1839);
   U9954 : OAI22_X1 port map( A1 => n10179, A2 => n9870, B1 => n7280, B2 => 
                           n9866, ZN => n1840);
   U9955 : OAI22_X1 port map( A1 => n10182, A2 => n9870, B1 => n7279, B2 => 
                           n9866, ZN => n1841);
   U9956 : OAI22_X1 port map( A1 => n10185, A2 => n9870, B1 => n7278, B2 => 
                           n9866, ZN => n1842);
   U9957 : OAI22_X1 port map( A1 => n10188, A2 => n9870, B1 => n7277, B2 => 
                           n9866, ZN => n1843);
   U9958 : OAI22_X1 port map( A1 => n10191, A2 => n9870, B1 => n7276, B2 => 
                           n9866, ZN => n1844);
   U9959 : OAI22_X1 port map( A1 => n10194, A2 => n9870, B1 => n7275, B2 => 
                           n9866, ZN => n1845);
   U9960 : OAI22_X1 port map( A1 => n10197, A2 => n9870, B1 => n7274, B2 => 
                           n9866, ZN => n1846);
   U9961 : OAI22_X1 port map( A1 => n10200, A2 => n9871, B1 => n7273, B2 => 
                           n9866, ZN => n1847);
   U9962 : OAI22_X1 port map( A1 => n10203, A2 => n9871, B1 => n7272, B2 => 
                           n9867, ZN => n1848);
   U9963 : OAI22_X1 port map( A1 => n10206, A2 => n9871, B1 => n7271, B2 => 
                           n9867, ZN => n1849);
   U9964 : OAI22_X1 port map( A1 => n10209, A2 => n9871, B1 => n7270, B2 => 
                           n9867, ZN => n1850);
   U9965 : OAI22_X1 port map( A1 => n10212, A2 => n9871, B1 => n7269, B2 => 
                           n9867, ZN => n1851);
   U9966 : OAI22_X1 port map( A1 => n10215, A2 => n9871, B1 => n7268, B2 => 
                           n9867, ZN => n1852);
   U9967 : OAI22_X1 port map( A1 => n10218, A2 => n9871, B1 => n7267, B2 => 
                           n9867, ZN => n1853);
   U9968 : OAI22_X1 port map( A1 => n10221, A2 => n9871, B1 => n7266, B2 => 
                           n9867, ZN => n1854);
   U9969 : OAI22_X1 port map( A1 => n10130, A2 => n9925, B1 => n7073, B2 => 
                           n9921, ZN => n2048);
   U9970 : OAI22_X1 port map( A1 => n10133, A2 => n9925, B1 => n7072, B2 => 
                           n9921, ZN => n2049);
   U9971 : OAI22_X1 port map( A1 => n10136, A2 => n9925, B1 => n7071, B2 => 
                           n9921, ZN => n2050);
   U9972 : OAI22_X1 port map( A1 => n10139, A2 => n9925, B1 => n7070, B2 => 
                           n9921, ZN => n2051);
   U9973 : OAI22_X1 port map( A1 => n10142, A2 => n9925, B1 => n7069, B2 => 
                           n9921, ZN => n2052);
   U9974 : OAI22_X1 port map( A1 => n10145, A2 => n9925, B1 => n7068, B2 => 
                           n9921, ZN => n2053);
   U9975 : OAI22_X1 port map( A1 => n10148, A2 => n9925, B1 => n7067, B2 => 
                           n9921, ZN => n2054);
   U9976 : OAI22_X1 port map( A1 => n10151, A2 => n9925, B1 => n7066, B2 => 
                           n9921, ZN => n2055);
   U9977 : OAI22_X1 port map( A1 => n10154, A2 => n9925, B1 => n7065, B2 => 
                           n9921, ZN => n2056);
   U9978 : OAI22_X1 port map( A1 => n10157, A2 => n9925, B1 => n7064, B2 => 
                           n9921, ZN => n2057);
   U9979 : OAI22_X1 port map( A1 => n10160, A2 => n9925, B1 => n7063, B2 => 
                           n9921, ZN => n2058);
   U9980 : OAI22_X1 port map( A1 => n10163, A2 => n9926, B1 => n7062, B2 => 
                           n9921, ZN => n2059);
   U9981 : OAI22_X1 port map( A1 => n10166, A2 => n9926, B1 => n7061, B2 => 
                           n9922, ZN => n2060);
   U9982 : OAI22_X1 port map( A1 => n10169, A2 => n9926, B1 => n7060, B2 => 
                           n9922, ZN => n2061);
   U9983 : OAI22_X1 port map( A1 => n10172, A2 => n9926, B1 => n7059, B2 => 
                           n9922, ZN => n2062);
   U9984 : OAI22_X1 port map( A1 => n10175, A2 => n9926, B1 => n7058, B2 => 
                           n9922, ZN => n2063);
   U9985 : OAI22_X1 port map( A1 => n10178, A2 => n9926, B1 => n7057, B2 => 
                           n9922, ZN => n2064);
   U9986 : OAI22_X1 port map( A1 => n10181, A2 => n9926, B1 => n7056, B2 => 
                           n9922, ZN => n2065);
   U9987 : OAI22_X1 port map( A1 => n10184, A2 => n9926, B1 => n7055, B2 => 
                           n9922, ZN => n2066);
   U9988 : OAI22_X1 port map( A1 => n10187, A2 => n9926, B1 => n7054, B2 => 
                           n9922, ZN => n2067);
   U9989 : OAI22_X1 port map( A1 => n10190, A2 => n9926, B1 => n7053, B2 => 
                           n9922, ZN => n2068);
   U9990 : OAI22_X1 port map( A1 => n10193, A2 => n9926, B1 => n7052, B2 => 
                           n9922, ZN => n2069);
   U9991 : OAI22_X1 port map( A1 => n10196, A2 => n9926, B1 => n7051, B2 => 
                           n9922, ZN => n2070);
   U9992 : OAI22_X1 port map( A1 => n10199, A2 => n9927, B1 => n7050, B2 => 
                           n9922, ZN => n2071);
   U9993 : OAI22_X1 port map( A1 => n10202, A2 => n9927, B1 => n7049, B2 => 
                           n9923, ZN => n2072);
   U9994 : OAI22_X1 port map( A1 => n10205, A2 => n9927, B1 => n7048, B2 => 
                           n9923, ZN => n2073);
   U9995 : OAI22_X1 port map( A1 => n10208, A2 => n9927, B1 => n7047, B2 => 
                           n9923, ZN => n2074);
   U9996 : OAI22_X1 port map( A1 => n10211, A2 => n9927, B1 => n7046, B2 => 
                           n9923, ZN => n2075);
   U9997 : OAI22_X1 port map( A1 => n10214, A2 => n9927, B1 => n7045, B2 => 
                           n9923, ZN => n2076);
   U9998 : OAI22_X1 port map( A1 => n10217, A2 => n9927, B1 => n7044, B2 => 
                           n9923, ZN => n2077);
   U9999 : OAI22_X1 port map( A1 => n10220, A2 => n9927, B1 => n7043, B2 => 
                           n9923, ZN => n2078);
   U10000 : OAI22_X1 port map( A1 => n10223, A2 => n9927, B1 => n7042, B2 => 
                           n9923, ZN => n2079);
   U10001 : OAI22_X1 port map( A1 => n10130, A2 => n9957, B1 => n6945, B2 => 
                           n9953, ZN => n2176);
   U10002 : OAI22_X1 port map( A1 => n10133, A2 => n9957, B1 => n6944, B2 => 
                           n9953, ZN => n2177);
   U10003 : OAI22_X1 port map( A1 => n10136, A2 => n9957, B1 => n6943, B2 => 
                           n9953, ZN => n2178);
   U10004 : OAI22_X1 port map( A1 => n10139, A2 => n9957, B1 => n6942, B2 => 
                           n9953, ZN => n2179);
   U10005 : OAI22_X1 port map( A1 => n10142, A2 => n9957, B1 => n6941, B2 => 
                           n9953, ZN => n2180);
   U10006 : OAI22_X1 port map( A1 => n10145, A2 => n9957, B1 => n6940, B2 => 
                           n9953, ZN => n2181);
   U10007 : OAI22_X1 port map( A1 => n10148, A2 => n9957, B1 => n6939, B2 => 
                           n9953, ZN => n2182);
   U10008 : OAI22_X1 port map( A1 => n10151, A2 => n9957, B1 => n6938, B2 => 
                           n9953, ZN => n2183);
   U10009 : OAI22_X1 port map( A1 => n10154, A2 => n9957, B1 => n6937, B2 => 
                           n9953, ZN => n2184);
   U10010 : OAI22_X1 port map( A1 => n10157, A2 => n9957, B1 => n6936, B2 => 
                           n9953, ZN => n2185);
   U10011 : OAI22_X1 port map( A1 => n10160, A2 => n9957, B1 => n6935, B2 => 
                           n9953, ZN => n2186);
   U10012 : OAI22_X1 port map( A1 => n10163, A2 => n9958, B1 => n6934, B2 => 
                           n9953, ZN => n2187);
   U10013 : OAI22_X1 port map( A1 => n10166, A2 => n9958, B1 => n6933, B2 => 
                           n9954, ZN => n2188);
   U10014 : OAI22_X1 port map( A1 => n10169, A2 => n9958, B1 => n6932, B2 => 
                           n9954, ZN => n2189);
   U10015 : OAI22_X1 port map( A1 => n10172, A2 => n9958, B1 => n6931, B2 => 
                           n9954, ZN => n2190);
   U10016 : OAI22_X1 port map( A1 => n10175, A2 => n9958, B1 => n6930, B2 => 
                           n9954, ZN => n2191);
   U10017 : OAI22_X1 port map( A1 => n10178, A2 => n9958, B1 => n6929, B2 => 
                           n9954, ZN => n2192);
   U10018 : OAI22_X1 port map( A1 => n10181, A2 => n9958, B1 => n6928, B2 => 
                           n9954, ZN => n2193);
   U10019 : OAI22_X1 port map( A1 => n10184, A2 => n9958, B1 => n6927, B2 => 
                           n9954, ZN => n2194);
   U10020 : OAI22_X1 port map( A1 => n10187, A2 => n9958, B1 => n6926, B2 => 
                           n9954, ZN => n2195);
   U10021 : OAI22_X1 port map( A1 => n10190, A2 => n9958, B1 => n6925, B2 => 
                           n9954, ZN => n2196);
   U10022 : OAI22_X1 port map( A1 => n10193, A2 => n9958, B1 => n6924, B2 => 
                           n9954, ZN => n2197);
   U10023 : OAI22_X1 port map( A1 => n10196, A2 => n9958, B1 => n6923, B2 => 
                           n9954, ZN => n2198);
   U10024 : OAI22_X1 port map( A1 => n10199, A2 => n9959, B1 => n6922, B2 => 
                           n9954, ZN => n2199);
   U10025 : OAI22_X1 port map( A1 => n10202, A2 => n9959, B1 => n6921, B2 => 
                           n9955, ZN => n2200);
   U10026 : OAI22_X1 port map( A1 => n10205, A2 => n9959, B1 => n6920, B2 => 
                           n9955, ZN => n2201);
   U10027 : OAI22_X1 port map( A1 => n10208, A2 => n9959, B1 => n6919, B2 => 
                           n9955, ZN => n2202);
   U10028 : OAI22_X1 port map( A1 => n10211, A2 => n9959, B1 => n6918, B2 => 
                           n9955, ZN => n2203);
   U10029 : OAI22_X1 port map( A1 => n10214, A2 => n9959, B1 => n6917, B2 => 
                           n9955, ZN => n2204);
   U10030 : OAI22_X1 port map( A1 => n10217, A2 => n9959, B1 => n6916, B2 => 
                           n9955, ZN => n2205);
   U10031 : OAI22_X1 port map( A1 => n10220, A2 => n9959, B1 => n6915, B2 => 
                           n9955, ZN => n2206);
   U10032 : OAI22_X1 port map( A1 => n10223, A2 => n9959, B1 => n6914, B2 => 
                           n9955, ZN => n2207);
   U10033 : OAI22_X1 port map( A1 => n10130, A2 => n9965, B1 => n6913, B2 => 
                           n9961, ZN => n2208);
   U10034 : OAI22_X1 port map( A1 => n10133, A2 => n9965, B1 => n6912, B2 => 
                           n9961, ZN => n2209);
   U10035 : OAI22_X1 port map( A1 => n10136, A2 => n9965, B1 => n6911, B2 => 
                           n9961, ZN => n2210);
   U10036 : OAI22_X1 port map( A1 => n10139, A2 => n9965, B1 => n6910, B2 => 
                           n9961, ZN => n2211);
   U10037 : OAI22_X1 port map( A1 => n10142, A2 => n9965, B1 => n6909, B2 => 
                           n9961, ZN => n2212);
   U10038 : OAI22_X1 port map( A1 => n10145, A2 => n9965, B1 => n6908, B2 => 
                           n9961, ZN => n2213);
   U10039 : OAI22_X1 port map( A1 => n10148, A2 => n9965, B1 => n6907, B2 => 
                           n9961, ZN => n2214);
   U10040 : OAI22_X1 port map( A1 => n10151, A2 => n9965, B1 => n6906, B2 => 
                           n9961, ZN => n2215);
   U10041 : OAI22_X1 port map( A1 => n10154, A2 => n9965, B1 => n6905, B2 => 
                           n9961, ZN => n2216);
   U10042 : OAI22_X1 port map( A1 => n10157, A2 => n9965, B1 => n6904, B2 => 
                           n9961, ZN => n2217);
   U10043 : OAI22_X1 port map( A1 => n10160, A2 => n9965, B1 => n6903, B2 => 
                           n9961, ZN => n2218);
   U10044 : OAI22_X1 port map( A1 => n10163, A2 => n9966, B1 => n6902, B2 => 
                           n9961, ZN => n2219);
   U10045 : OAI22_X1 port map( A1 => n10166, A2 => n9966, B1 => n6901, B2 => 
                           n9962, ZN => n2220);
   U10046 : OAI22_X1 port map( A1 => n10169, A2 => n9966, B1 => n6900, B2 => 
                           n9962, ZN => n2221);
   U10047 : OAI22_X1 port map( A1 => n10172, A2 => n9966, B1 => n6899, B2 => 
                           n9962, ZN => n2222);
   U10048 : OAI22_X1 port map( A1 => n10175, A2 => n9966, B1 => n6898, B2 => 
                           n9962, ZN => n2223);
   U10049 : OAI22_X1 port map( A1 => n10178, A2 => n9966, B1 => n6897, B2 => 
                           n9962, ZN => n2224);
   U10050 : OAI22_X1 port map( A1 => n10181, A2 => n9966, B1 => n6896, B2 => 
                           n9962, ZN => n2225);
   U10051 : OAI22_X1 port map( A1 => n10184, A2 => n9966, B1 => n6895, B2 => 
                           n9962, ZN => n2226);
   U10052 : OAI22_X1 port map( A1 => n10187, A2 => n9966, B1 => n6894, B2 => 
                           n9962, ZN => n2227);
   U10053 : OAI22_X1 port map( A1 => n10190, A2 => n9966, B1 => n6893, B2 => 
                           n9962, ZN => n2228);
   U10054 : OAI22_X1 port map( A1 => n10193, A2 => n9966, B1 => n6892, B2 => 
                           n9962, ZN => n2229);
   U10055 : OAI22_X1 port map( A1 => n10196, A2 => n9966, B1 => n6891, B2 => 
                           n9962, ZN => n2230);
   U10056 : OAI22_X1 port map( A1 => n10199, A2 => n9967, B1 => n6890, B2 => 
                           n9962, ZN => n2231);
   U10057 : OAI22_X1 port map( A1 => n10202, A2 => n9967, B1 => n6889, B2 => 
                           n9963, ZN => n2232);
   U10058 : OAI22_X1 port map( A1 => n10205, A2 => n9967, B1 => n6888, B2 => 
                           n9963, ZN => n2233);
   U10059 : OAI22_X1 port map( A1 => n10208, A2 => n9967, B1 => n6887, B2 => 
                           n9963, ZN => n2234);
   U10060 : OAI22_X1 port map( A1 => n10211, A2 => n9967, B1 => n6886, B2 => 
                           n9963, ZN => n2235);
   U10061 : OAI22_X1 port map( A1 => n10214, A2 => n9967, B1 => n6885, B2 => 
                           n9963, ZN => n2236);
   U10062 : OAI22_X1 port map( A1 => n10217, A2 => n9967, B1 => n6884, B2 => 
                           n9963, ZN => n2237);
   U10063 : OAI22_X1 port map( A1 => n10220, A2 => n9967, B1 => n6883, B2 => 
                           n9963, ZN => n2238);
   U10064 : OAI22_X1 port map( A1 => n10223, A2 => n9967, B1 => n6882, B2 => 
                           n9963, ZN => n2239);
   U10065 : OAI22_X1 port map( A1 => n10131, A2 => n9861, B1 => n704, B2 => 
                           n9857, ZN => n1792);
   U10066 : OAI22_X1 port map( A1 => n10134, A2 => n9861, B1 => n705, B2 => 
                           n9857, ZN => n1793);
   U10067 : OAI22_X1 port map( A1 => n10137, A2 => n9861, B1 => n706, B2 => 
                           n9857, ZN => n1794);
   U10068 : OAI22_X1 port map( A1 => n10140, A2 => n9861, B1 => n707, B2 => 
                           n9857, ZN => n1795);
   U10069 : OAI22_X1 port map( A1 => n10143, A2 => n9861, B1 => n708, B2 => 
                           n9857, ZN => n1796);
   U10070 : OAI22_X1 port map( A1 => n10146, A2 => n9861, B1 => n709, B2 => 
                           n9857, ZN => n1797);
   U10071 : OAI22_X1 port map( A1 => n10149, A2 => n9861, B1 => n710, B2 => 
                           n9857, ZN => n1798);
   U10072 : OAI22_X1 port map( A1 => n10152, A2 => n9861, B1 => n711, B2 => 
                           n9857, ZN => n1799);
   U10073 : OAI22_X1 port map( A1 => n10155, A2 => n9861, B1 => n712, B2 => 
                           n9857, ZN => n1800);
   U10074 : OAI22_X1 port map( A1 => n10158, A2 => n9861, B1 => n713, B2 => 
                           n9857, ZN => n1801);
   U10075 : OAI22_X1 port map( A1 => n10161, A2 => n9861, B1 => n714, B2 => 
                           n9857, ZN => n1802);
   U10076 : OAI22_X1 port map( A1 => n10164, A2 => n9862, B1 => n715, B2 => 
                           n9857, ZN => n1803);
   U10077 : OAI22_X1 port map( A1 => n10167, A2 => n9862, B1 => n716, B2 => 
                           n9858, ZN => n1804);
   U10078 : OAI22_X1 port map( A1 => n10170, A2 => n9862, B1 => n717, B2 => 
                           n9858, ZN => n1805);
   U10079 : OAI22_X1 port map( A1 => n10173, A2 => n9862, B1 => n718, B2 => 
                           n9858, ZN => n1806);
   U10080 : OAI22_X1 port map( A1 => n10176, A2 => n9862, B1 => n719, B2 => 
                           n9858, ZN => n1807);
   U10081 : OAI22_X1 port map( A1 => n10179, A2 => n9862, B1 => n720, B2 => 
                           n9858, ZN => n1808);
   U10082 : OAI22_X1 port map( A1 => n10182, A2 => n9862, B1 => n721, B2 => 
                           n9858, ZN => n1809);
   U10083 : OAI22_X1 port map( A1 => n10185, A2 => n9862, B1 => n722, B2 => 
                           n9858, ZN => n1810);
   U10084 : OAI22_X1 port map( A1 => n10188, A2 => n9862, B1 => n723, B2 => 
                           n9858, ZN => n1811);
   U10085 : OAI22_X1 port map( A1 => n10191, A2 => n9862, B1 => n724, B2 => 
                           n9858, ZN => n1812);
   U10086 : OAI22_X1 port map( A1 => n10194, A2 => n9862, B1 => n725, B2 => 
                           n9858, ZN => n1813);
   U10087 : OAI22_X1 port map( A1 => n10197, A2 => n9862, B1 => n726, B2 => 
                           n9858, ZN => n1814);
   U10088 : OAI22_X1 port map( A1 => n10200, A2 => n9863, B1 => n727, B2 => 
                           n9858, ZN => n1815);
   U10089 : OAI22_X1 port map( A1 => n10131, A2 => n9845, B1 => n640, B2 => 
                           n9841, ZN => n1728);
   U10090 : OAI22_X1 port map( A1 => n10134, A2 => n9845, B1 => n641, B2 => 
                           n9841, ZN => n1729);
   U10091 : OAI22_X1 port map( A1 => n10137, A2 => n9845, B1 => n642, B2 => 
                           n9841, ZN => n1730);
   U10092 : OAI22_X1 port map( A1 => n10140, A2 => n9845, B1 => n643, B2 => 
                           n9841, ZN => n1731);
   U10093 : OAI22_X1 port map( A1 => n10143, A2 => n9845, B1 => n644, B2 => 
                           n9841, ZN => n1732);
   U10094 : OAI22_X1 port map( A1 => n10146, A2 => n9845, B1 => n645, B2 => 
                           n9841, ZN => n1733);
   U10095 : OAI22_X1 port map( A1 => n10149, A2 => n9845, B1 => n646, B2 => 
                           n9841, ZN => n1734);
   U10096 : OAI22_X1 port map( A1 => n10152, A2 => n9845, B1 => n647, B2 => 
                           n9841, ZN => n1735);
   U10097 : OAI22_X1 port map( A1 => n10155, A2 => n9845, B1 => n648, B2 => 
                           n9841, ZN => n1736);
   U10098 : OAI22_X1 port map( A1 => n10158, A2 => n9845, B1 => n649, B2 => 
                           n9841, ZN => n1737);
   U10099 : OAI22_X1 port map( A1 => n10161, A2 => n9845, B1 => n650, B2 => 
                           n9841, ZN => n1738);
   U10100 : OAI22_X1 port map( A1 => n10164, A2 => n9846, B1 => n651, B2 => 
                           n9841, ZN => n1739);
   U10101 : OAI22_X1 port map( A1 => n10167, A2 => n9846, B1 => n652, B2 => 
                           n9842, ZN => n1740);
   U10102 : OAI22_X1 port map( A1 => n10170, A2 => n9846, B1 => n653, B2 => 
                           n9842, ZN => n1741);
   U10103 : OAI22_X1 port map( A1 => n10173, A2 => n9846, B1 => n654, B2 => 
                           n9842, ZN => n1742);
   U10104 : OAI22_X1 port map( A1 => n10176, A2 => n9846, B1 => n655, B2 => 
                           n9842, ZN => n1743);
   U10105 : OAI22_X1 port map( A1 => n10179, A2 => n9846, B1 => n656, B2 => 
                           n9842, ZN => n1744);
   U10106 : OAI22_X1 port map( A1 => n10182, A2 => n9846, B1 => n657, B2 => 
                           n9842, ZN => n1745);
   U10107 : OAI22_X1 port map( A1 => n10185, A2 => n9846, B1 => n658, B2 => 
                           n9842, ZN => n1746);
   U10108 : OAI22_X1 port map( A1 => n10188, A2 => n9846, B1 => n659, B2 => 
                           n9842, ZN => n1747);
   U10109 : OAI22_X1 port map( A1 => n10191, A2 => n9846, B1 => n660, B2 => 
                           n9842, ZN => n1748);
   U10110 : OAI22_X1 port map( A1 => n10194, A2 => n9846, B1 => n661, B2 => 
                           n9842, ZN => n1749);
   U10111 : OAI22_X1 port map( A1 => n10197, A2 => n9846, B1 => n662, B2 => 
                           n9842, ZN => n1750);
   U10112 : OAI22_X1 port map( A1 => n10200, A2 => n9847, B1 => n663, B2 => 
                           n9842, ZN => n1751);
   U10113 : OAI22_X1 port map( A1 => n10131, A2 => n9805, B1 => n480, B2 => 
                           n9801, ZN => n1568);
   U10114 : OAI22_X1 port map( A1 => n10134, A2 => n9805, B1 => n481, B2 => 
                           n9801, ZN => n1569);
   U10115 : OAI22_X1 port map( A1 => n10137, A2 => n9805, B1 => n482, B2 => 
                           n9801, ZN => n1570);
   U10116 : OAI22_X1 port map( A1 => n10140, A2 => n9805, B1 => n483, B2 => 
                           n9801, ZN => n1571);
   U10117 : OAI22_X1 port map( A1 => n10143, A2 => n9805, B1 => n484, B2 => 
                           n9801, ZN => n1572);
   U10118 : OAI22_X1 port map( A1 => n10146, A2 => n9805, B1 => n485, B2 => 
                           n9801, ZN => n1573);
   U10119 : OAI22_X1 port map( A1 => n10149, A2 => n9805, B1 => n486, B2 => 
                           n9801, ZN => n1574);
   U10120 : OAI22_X1 port map( A1 => n10152, A2 => n9805, B1 => n487, B2 => 
                           n9801, ZN => n1575);
   U10121 : OAI22_X1 port map( A1 => n10155, A2 => n9805, B1 => n488, B2 => 
                           n9801, ZN => n1576);
   U10122 : OAI22_X1 port map( A1 => n10158, A2 => n9805, B1 => n489, B2 => 
                           n9801, ZN => n1577);
   U10123 : OAI22_X1 port map( A1 => n10161, A2 => n9805, B1 => n490, B2 => 
                           n9801, ZN => n1578);
   U10124 : OAI22_X1 port map( A1 => n10164, A2 => n9806, B1 => n491, B2 => 
                           n9801, ZN => n1579);
   U10125 : OAI22_X1 port map( A1 => n10167, A2 => n9806, B1 => n492, B2 => 
                           n9802, ZN => n1580);
   U10126 : OAI22_X1 port map( A1 => n10170, A2 => n9806, B1 => n493, B2 => 
                           n9802, ZN => n1581);
   U10127 : OAI22_X1 port map( A1 => n10173, A2 => n9806, B1 => n494, B2 => 
                           n9802, ZN => n1582);
   U10128 : OAI22_X1 port map( A1 => n10176, A2 => n9806, B1 => n495, B2 => 
                           n9802, ZN => n1583);
   U10129 : OAI22_X1 port map( A1 => n10179, A2 => n9806, B1 => n496, B2 => 
                           n9802, ZN => n1584);
   U10130 : OAI22_X1 port map( A1 => n10182, A2 => n9806, B1 => n497, B2 => 
                           n9802, ZN => n1585);
   U10131 : OAI22_X1 port map( A1 => n10185, A2 => n9806, B1 => n498, B2 => 
                           n9802, ZN => n1586);
   U10132 : OAI22_X1 port map( A1 => n10188, A2 => n9806, B1 => n499, B2 => 
                           n9802, ZN => n1587);
   U10133 : OAI22_X1 port map( A1 => n10191, A2 => n9806, B1 => n500, B2 => 
                           n9802, ZN => n1588);
   U10134 : OAI22_X1 port map( A1 => n10194, A2 => n9806, B1 => n501, B2 => 
                           n9802, ZN => n1589);
   U10135 : OAI22_X1 port map( A1 => n10197, A2 => n9806, B1 => n502, B2 => 
                           n9802, ZN => n1590);
   U10136 : OAI22_X1 port map( A1 => n10200, A2 => n9807, B1 => n503, B2 => 
                           n9802, ZN => n1591);
   U10137 : OAI22_X1 port map( A1 => n10179, A2 => n9798, B1 => n464, B2 => 
                           n9794, ZN => n1552);
   U10138 : OAI22_X1 port map( A1 => n10182, A2 => n9798, B1 => n465, B2 => 
                           n9794, ZN => n1553);
   U10139 : OAI22_X1 port map( A1 => n10185, A2 => n9798, B1 => n466, B2 => 
                           n9794, ZN => n1554);
   U10140 : OAI22_X1 port map( A1 => n10188, A2 => n9798, B1 => n467, B2 => 
                           n9794, ZN => n1555);
   U10141 : OAI22_X1 port map( A1 => n10191, A2 => n9798, B1 => n468, B2 => 
                           n9794, ZN => n1556);
   U10142 : OAI22_X1 port map( A1 => n10194, A2 => n9798, B1 => n469, B2 => 
                           n9794, ZN => n1557);
   U10143 : OAI22_X1 port map( A1 => n10197, A2 => n9798, B1 => n470, B2 => 
                           n9794, ZN => n1558);
   U10144 : OAI22_X1 port map( A1 => n10200, A2 => n9799, B1 => n471, B2 => 
                           n9794, ZN => n1559);
   U10145 : OAI22_X1 port map( A1 => n10203, A2 => n9863, B1 => n728, B2 => 
                           n9859, ZN => n1816);
   U10146 : OAI22_X1 port map( A1 => n10206, A2 => n9863, B1 => n729, B2 => 
                           n9859, ZN => n1817);
   U10147 : OAI22_X1 port map( A1 => n10209, A2 => n9863, B1 => n730, B2 => 
                           n9859, ZN => n1818);
   U10148 : OAI22_X1 port map( A1 => n10212, A2 => n9863, B1 => n731, B2 => 
                           n9859, ZN => n1819);
   U10149 : OAI22_X1 port map( A1 => n10215, A2 => n9863, B1 => n732, B2 => 
                           n9859, ZN => n1820);
   U10150 : OAI22_X1 port map( A1 => n10218, A2 => n9863, B1 => n733, B2 => 
                           n9859, ZN => n1821);
   U10151 : OAI22_X1 port map( A1 => n10221, A2 => n9863, B1 => n734, B2 => 
                           n9859, ZN => n1822);
   U10152 : OAI22_X1 port map( A1 => n10224, A2 => n9863, B1 => n735, B2 => 
                           n9859, ZN => n1823);
   U10153 : OAI22_X1 port map( A1 => n10203, A2 => n9847, B1 => n664, B2 => 
                           n9843, ZN => n1752);
   U10154 : OAI22_X1 port map( A1 => n10206, A2 => n9847, B1 => n665, B2 => 
                           n9843, ZN => n1753);
   U10155 : OAI22_X1 port map( A1 => n10209, A2 => n9847, B1 => n666, B2 => 
                           n9843, ZN => n1754);
   U10156 : OAI22_X1 port map( A1 => n10212, A2 => n9847, B1 => n667, B2 => 
                           n9843, ZN => n1755);
   U10157 : OAI22_X1 port map( A1 => n10215, A2 => n9847, B1 => n668, B2 => 
                           n9843, ZN => n1756);
   U10158 : OAI22_X1 port map( A1 => n10218, A2 => n9847, B1 => n669, B2 => 
                           n9843, ZN => n1757);
   U10159 : OAI22_X1 port map( A1 => n10221, A2 => n9847, B1 => n670, B2 => 
                           n9843, ZN => n1758);
   U10160 : OAI22_X1 port map( A1 => n10224, A2 => n9847, B1 => n671, B2 => 
                           n9843, ZN => n1759);
   U10161 : OAI22_X1 port map( A1 => n10203, A2 => n9807, B1 => n504, B2 => 
                           n9803, ZN => n1592);
   U10162 : OAI22_X1 port map( A1 => n10206, A2 => n9807, B1 => n505, B2 => 
                           n9803, ZN => n1593);
   U10163 : OAI22_X1 port map( A1 => n10209, A2 => n9807, B1 => n506, B2 => 
                           n9803, ZN => n1594);
   U10164 : OAI22_X1 port map( A1 => n10212, A2 => n9807, B1 => n507, B2 => 
                           n9803, ZN => n1595);
   U10165 : OAI22_X1 port map( A1 => n10215, A2 => n9807, B1 => n508, B2 => 
                           n9803, ZN => n1596);
   U10166 : OAI22_X1 port map( A1 => n10218, A2 => n9807, B1 => n509, B2 => 
                           n9803, ZN => n1597);
   U10167 : OAI22_X1 port map( A1 => n10221, A2 => n9807, B1 => n510, B2 => 
                           n9803, ZN => n1598);
   U10168 : OAI22_X1 port map( A1 => n10224, A2 => n9807, B1 => n511, B2 => 
                           n9803, ZN => n1599);
   U10169 : OAI22_X1 port map( A1 => n10203, A2 => n9799, B1 => n472, B2 => 
                           n9795, ZN => n1560);
   U10170 : OAI22_X1 port map( A1 => n10206, A2 => n9799, B1 => n473, B2 => 
                           n9795, ZN => n1561);
   U10171 : OAI22_X1 port map( A1 => n10209, A2 => n9799, B1 => n474, B2 => 
                           n9795, ZN => n1562);
   U10172 : OAI22_X1 port map( A1 => n10212, A2 => n9799, B1 => n475, B2 => 
                           n9795, ZN => n1563);
   U10173 : OAI22_X1 port map( A1 => n10215, A2 => n9799, B1 => n476, B2 => 
                           n9795, ZN => n1564);
   U10174 : OAI22_X1 port map( A1 => n10218, A2 => n9799, B1 => n477, B2 => 
                           n9795, ZN => n1565);
   U10175 : OAI22_X1 port map( A1 => n10221, A2 => n9799, B1 => n478, B2 => 
                           n9795, ZN => n1566);
   U10176 : OAI22_X1 port map( A1 => n10224, A2 => n9799, B1 => n479, B2 => 
                           n9795, ZN => n1567);
   U10177 : OAI22_X1 port map( A1 => n10131, A2 => n9821, B1 => n544, B2 => 
                           n9817, ZN => n1632);
   U10178 : OAI22_X1 port map( A1 => n10134, A2 => n9821, B1 => n545, B2 => 
                           n9817, ZN => n1633);
   U10179 : OAI22_X1 port map( A1 => n10137, A2 => n9821, B1 => n546, B2 => 
                           n9817, ZN => n1634);
   U10180 : OAI22_X1 port map( A1 => n10140, A2 => n9821, B1 => n547, B2 => 
                           n9817, ZN => n1635);
   U10181 : OAI22_X1 port map( A1 => n10143, A2 => n9821, B1 => n548, B2 => 
                           n9817, ZN => n1636);
   U10182 : OAI22_X1 port map( A1 => n10146, A2 => n9821, B1 => n549, B2 => 
                           n9817, ZN => n1637);
   U10183 : OAI22_X1 port map( A1 => n10149, A2 => n9821, B1 => n550, B2 => 
                           n9817, ZN => n1638);
   U10184 : OAI22_X1 port map( A1 => n10152, A2 => n9821, B1 => n551, B2 => 
                           n9817, ZN => n1639);
   U10185 : OAI22_X1 port map( A1 => n10155, A2 => n9821, B1 => n552, B2 => 
                           n9817, ZN => n1640);
   U10186 : OAI22_X1 port map( A1 => n10158, A2 => n9821, B1 => n553, B2 => 
                           n9817, ZN => n1641);
   U10187 : OAI22_X1 port map( A1 => n10161, A2 => n9821, B1 => n554, B2 => 
                           n9817, ZN => n1642);
   U10188 : OAI22_X1 port map( A1 => n10164, A2 => n9822, B1 => n555, B2 => 
                           n9817, ZN => n1643);
   U10189 : OAI22_X1 port map( A1 => n10167, A2 => n9822, B1 => n556, B2 => 
                           n9818, ZN => n1644);
   U10190 : OAI22_X1 port map( A1 => n10170, A2 => n9822, B1 => n557, B2 => 
                           n9818, ZN => n1645);
   U10191 : OAI22_X1 port map( A1 => n10173, A2 => n9822, B1 => n558, B2 => 
                           n9818, ZN => n1646);
   U10192 : OAI22_X1 port map( A1 => n10176, A2 => n9822, B1 => n559, B2 => 
                           n9818, ZN => n1647);
   U10193 : OAI22_X1 port map( A1 => n10179, A2 => n9822, B1 => n560, B2 => 
                           n9818, ZN => n1648);
   U10194 : OAI22_X1 port map( A1 => n10182, A2 => n9822, B1 => n561, B2 => 
                           n9818, ZN => n1649);
   U10195 : OAI22_X1 port map( A1 => n10185, A2 => n9822, B1 => n562, B2 => 
                           n9818, ZN => n1650);
   U10196 : OAI22_X1 port map( A1 => n10188, A2 => n9822, B1 => n563, B2 => 
                           n9818, ZN => n1651);
   U10197 : OAI22_X1 port map( A1 => n10191, A2 => n9822, B1 => n564, B2 => 
                           n9818, ZN => n1652);
   U10198 : OAI22_X1 port map( A1 => n10194, A2 => n9822, B1 => n565, B2 => 
                           n9818, ZN => n1653);
   U10199 : OAI22_X1 port map( A1 => n10197, A2 => n9822, B1 => n566, B2 => 
                           n9818, ZN => n1654);
   U10200 : OAI22_X1 port map( A1 => n10200, A2 => n9823, B1 => n567, B2 => 
                           n9818, ZN => n1655);
   U10201 : OAI22_X1 port map( A1 => n10131, A2 => n9813, B1 => n512, B2 => 
                           n9809, ZN => n1600);
   U10202 : OAI22_X1 port map( A1 => n10134, A2 => n9813, B1 => n513, B2 => 
                           n9809, ZN => n1601);
   U10203 : OAI22_X1 port map( A1 => n10137, A2 => n9813, B1 => n514, B2 => 
                           n9809, ZN => n1602);
   U10204 : OAI22_X1 port map( A1 => n10140, A2 => n9813, B1 => n515, B2 => 
                           n9809, ZN => n1603);
   U10205 : OAI22_X1 port map( A1 => n10143, A2 => n9813, B1 => n516, B2 => 
                           n9809, ZN => n1604);
   U10206 : OAI22_X1 port map( A1 => n10146, A2 => n9813, B1 => n517, B2 => 
                           n9809, ZN => n1605);
   U10207 : OAI22_X1 port map( A1 => n10149, A2 => n9813, B1 => n518, B2 => 
                           n9809, ZN => n1606);
   U10208 : OAI22_X1 port map( A1 => n10152, A2 => n9813, B1 => n519, B2 => 
                           n9809, ZN => n1607);
   U10209 : OAI22_X1 port map( A1 => n10155, A2 => n9813, B1 => n520, B2 => 
                           n9809, ZN => n1608);
   U10210 : OAI22_X1 port map( A1 => n10158, A2 => n9813, B1 => n521, B2 => 
                           n9809, ZN => n1609);
   U10211 : OAI22_X1 port map( A1 => n10161, A2 => n9813, B1 => n522, B2 => 
                           n9809, ZN => n1610);
   U10212 : OAI22_X1 port map( A1 => n10164, A2 => n9814, B1 => n523, B2 => 
                           n9809, ZN => n1611);
   U10213 : OAI22_X1 port map( A1 => n10167, A2 => n9814, B1 => n524, B2 => 
                           n9810, ZN => n1612);
   U10214 : OAI22_X1 port map( A1 => n10170, A2 => n9814, B1 => n525, B2 => 
                           n9810, ZN => n1613);
   U10215 : OAI22_X1 port map( A1 => n10173, A2 => n9814, B1 => n526, B2 => 
                           n9810, ZN => n1614);
   U10216 : OAI22_X1 port map( A1 => n10176, A2 => n9814, B1 => n527, B2 => 
                           n9810, ZN => n1615);
   U10217 : OAI22_X1 port map( A1 => n10179, A2 => n9814, B1 => n528, B2 => 
                           n9810, ZN => n1616);
   U10218 : OAI22_X1 port map( A1 => n10182, A2 => n9814, B1 => n529, B2 => 
                           n9810, ZN => n1617);
   U10219 : OAI22_X1 port map( A1 => n10185, A2 => n9814, B1 => n530, B2 => 
                           n9810, ZN => n1618);
   U10220 : OAI22_X1 port map( A1 => n10188, A2 => n9814, B1 => n531, B2 => 
                           n9810, ZN => n1619);
   U10221 : OAI22_X1 port map( A1 => n10191, A2 => n9814, B1 => n532, B2 => 
                           n9810, ZN => n1620);
   U10222 : OAI22_X1 port map( A1 => n10194, A2 => n9814, B1 => n533, B2 => 
                           n9810, ZN => n1621);
   U10223 : OAI22_X1 port map( A1 => n10197, A2 => n9814, B1 => n534, B2 => 
                           n9810, ZN => n1622);
   U10224 : OAI22_X1 port map( A1 => n10200, A2 => n9815, B1 => n535, B2 => 
                           n9810, ZN => n1623);
   U10225 : OAI22_X1 port map( A1 => n10203, A2 => n9823, B1 => n568, B2 => 
                           n9819, ZN => n1656);
   U10226 : OAI22_X1 port map( A1 => n10206, A2 => n9823, B1 => n569, B2 => 
                           n9819, ZN => n1657);
   U10227 : OAI22_X1 port map( A1 => n10209, A2 => n9823, B1 => n570, B2 => 
                           n9819, ZN => n1658);
   U10228 : OAI22_X1 port map( A1 => n10212, A2 => n9823, B1 => n571, B2 => 
                           n9819, ZN => n1659);
   U10229 : OAI22_X1 port map( A1 => n10215, A2 => n9823, B1 => n572, B2 => 
                           n9819, ZN => n1660);
   U10230 : OAI22_X1 port map( A1 => n10218, A2 => n9823, B1 => n573, B2 => 
                           n9819, ZN => n1661);
   U10231 : OAI22_X1 port map( A1 => n10221, A2 => n9823, B1 => n574, B2 => 
                           n9819, ZN => n1662);
   U10232 : OAI22_X1 port map( A1 => n10224, A2 => n9823, B1 => n575, B2 => 
                           n9819, ZN => n1663);
   U10233 : OAI22_X1 port map( A1 => n10203, A2 => n9815, B1 => n536, B2 => 
                           n9811, ZN => n1624);
   U10234 : OAI22_X1 port map( A1 => n10206, A2 => n9815, B1 => n537, B2 => 
                           n9811, ZN => n1625);
   U10235 : OAI22_X1 port map( A1 => n10209, A2 => n9815, B1 => n538, B2 => 
                           n9811, ZN => n1626);
   U10236 : OAI22_X1 port map( A1 => n10212, A2 => n9815, B1 => n539, B2 => 
                           n9811, ZN => n1627);
   U10237 : OAI22_X1 port map( A1 => n10215, A2 => n9815, B1 => n540, B2 => 
                           n9811, ZN => n1628);
   U10238 : OAI22_X1 port map( A1 => n10218, A2 => n9815, B1 => n541, B2 => 
                           n9811, ZN => n1629);
   U10239 : OAI22_X1 port map( A1 => n10221, A2 => n9815, B1 => n542, B2 => 
                           n9811, ZN => n1630);
   U10240 : OAI22_X1 port map( A1 => n10224, A2 => n9815, B1 => n543, B2 => 
                           n9811, ZN => n1631);
   U10241 : OAI22_X1 port map( A1 => n10131, A2 => n9829, B1 => n576, B2 => 
                           n9825, ZN => n1664);
   U10242 : OAI22_X1 port map( A1 => n10134, A2 => n9829, B1 => n577, B2 => 
                           n9825, ZN => n1665);
   U10243 : OAI22_X1 port map( A1 => n10137, A2 => n9829, B1 => n578, B2 => 
                           n9825, ZN => n1666);
   U10244 : OAI22_X1 port map( A1 => n10140, A2 => n9829, B1 => n579, B2 => 
                           n9825, ZN => n1667);
   U10245 : OAI22_X1 port map( A1 => n10143, A2 => n9829, B1 => n580, B2 => 
                           n9825, ZN => n1668);
   U10246 : OAI22_X1 port map( A1 => n10146, A2 => n9829, B1 => n581, B2 => 
                           n9825, ZN => n1669);
   U10247 : OAI22_X1 port map( A1 => n10149, A2 => n9829, B1 => n582, B2 => 
                           n9825, ZN => n1670);
   U10248 : OAI22_X1 port map( A1 => n10152, A2 => n9829, B1 => n583, B2 => 
                           n9825, ZN => n1671);
   U10249 : OAI22_X1 port map( A1 => n10155, A2 => n9829, B1 => n584, B2 => 
                           n9825, ZN => n1672);
   U10250 : OAI22_X1 port map( A1 => n10158, A2 => n9829, B1 => n585, B2 => 
                           n9825, ZN => n1673);
   U10251 : OAI22_X1 port map( A1 => n10161, A2 => n9829, B1 => n586, B2 => 
                           n9825, ZN => n1674);
   U10252 : OAI22_X1 port map( A1 => n10164, A2 => n9830, B1 => n587, B2 => 
                           n9825, ZN => n1675);
   U10253 : OAI22_X1 port map( A1 => n10167, A2 => n9830, B1 => n588, B2 => 
                           n9826, ZN => n1676);
   U10254 : OAI22_X1 port map( A1 => n10170, A2 => n9830, B1 => n589, B2 => 
                           n9826, ZN => n1677);
   U10255 : OAI22_X1 port map( A1 => n10173, A2 => n9830, B1 => n590, B2 => 
                           n9826, ZN => n1678);
   U10256 : OAI22_X1 port map( A1 => n10176, A2 => n9830, B1 => n591, B2 => 
                           n9826, ZN => n1679);
   U10257 : OAI22_X1 port map( A1 => n10179, A2 => n9830, B1 => n592, B2 => 
                           n9826, ZN => n1680);
   U10258 : OAI22_X1 port map( A1 => n10182, A2 => n9830, B1 => n593, B2 => 
                           n9826, ZN => n1681);
   U10259 : OAI22_X1 port map( A1 => n10185, A2 => n9830, B1 => n594, B2 => 
                           n9826, ZN => n1682);
   U10260 : OAI22_X1 port map( A1 => n10188, A2 => n9830, B1 => n595, B2 => 
                           n9826, ZN => n1683);
   U10261 : OAI22_X1 port map( A1 => n10191, A2 => n9830, B1 => n596, B2 => 
                           n9826, ZN => n1684);
   U10262 : OAI22_X1 port map( A1 => n10194, A2 => n9830, B1 => n597, B2 => 
                           n9826, ZN => n1685);
   U10263 : OAI22_X1 port map( A1 => n10197, A2 => n9830, B1 => n598, B2 => 
                           n9826, ZN => n1686);
   U10264 : OAI22_X1 port map( A1 => n10200, A2 => n9831, B1 => n599, B2 => 
                           n9826, ZN => n1687);
   U10265 : OAI22_X1 port map( A1 => n10203, A2 => n9831, B1 => n600, B2 => 
                           n9827, ZN => n1688);
   U10266 : OAI22_X1 port map( A1 => n10206, A2 => n9831, B1 => n601, B2 => 
                           n9827, ZN => n1689);
   U10267 : OAI22_X1 port map( A1 => n10209, A2 => n9831, B1 => n602, B2 => 
                           n9827, ZN => n1690);
   U10268 : OAI22_X1 port map( A1 => n10212, A2 => n9831, B1 => n603, B2 => 
                           n9827, ZN => n1691);
   U10269 : OAI22_X1 port map( A1 => n10215, A2 => n9831, B1 => n604, B2 => 
                           n9827, ZN => n1692);
   U10270 : OAI22_X1 port map( A1 => n10218, A2 => n9831, B1 => n605, B2 => 
                           n9827, ZN => n1693);
   U10271 : OAI22_X1 port map( A1 => n10221, A2 => n9831, B1 => n606, B2 => 
                           n9827, ZN => n1694);
   U10272 : OAI22_X1 port map( A1 => n10224, A2 => n9831, B1 => n607, B2 => 
                           n9827, ZN => n1695);
   U10273 : NOR3_X1 port map( A1 => n6747, A2 => ADD_RD1(1), A3 => n6749, ZN =>
                           n8878);
   U10274 : NOR3_X1 port map( A1 => n6751, A2 => ADD_RD2(1), A3 => n6753, ZN =>
                           n8210);
   U10275 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n8887);
   U10276 : NOR2_X1 port map( A1 => n6746, A2 => ADD_RD1(4), ZN => n8888);
   U10277 : NOR2_X1 port map( A1 => n6750, A2 => ADD_RD2(4), ZN => n8220);
   U10278 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n8219);
   U10279 : NOR3_X1 port map( A1 => n6748, A2 => ADD_RD1(0), A3 => n6747, ZN =>
                           n8869);
   U10280 : NOR3_X1 port map( A1 => n6752, A2 => ADD_RD2(0), A3 => n6751, ZN =>
                           n8201);
   U10281 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n6749, 
                           ZN => n8871);
   U10282 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n6753, 
                           ZN => n8203);
   U10283 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n6748, 
                           ZN => n8875);
   U10284 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n6752, 
                           ZN => n8207);
   U10285 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n8870);
   U10286 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n8202);
   U10287 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n6747, 
                           ZN => n8872);
   U10288 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n6751, 
                           ZN => n8204);
   U10289 : NOR3_X1 port map( A1 => n6748, A2 => ADD_RD1(2), A3 => n6749, ZN =>
                           n8874);
   U10290 : NOR3_X1 port map( A1 => n6752, A2 => ADD_RD2(2), A3 => n6753, ZN =>
                           n8206);
   U10291 : AND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n8236);
   U10292 : AND2_X1 port map( A1 => ADD_WR(1), A2 => n6745, ZN => n8233);
   U10293 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n6746, ZN => n8868);
   U10294 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n6750, ZN => n8200);
   U10295 : AND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n8876);
   U10296 : AND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n8208);
   U10297 : AND3_X1 port map( A1 => ADD_WR(2), A2 => n6743, A3 => n8274, ZN => 
                           n8277);
   U10298 : AND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n8274, ZN
                           => n8295);
   U10299 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n6744, A3 => n8274, ZN => 
                           n8286);
   U10300 : AND3_X1 port map( A1 => ADD_WR(2), A2 => n8237, A3 => ADD_WR(3), ZN
                           => n8258);
   U10301 : AND3_X1 port map( A1 => n8237, A2 => n6744, A3 => ADD_WR(3), ZN => 
                           n8249);
   U10302 : AND3_X1 port map( A1 => n8237, A2 => n6743, A3 => ADD_WR(2), ZN => 
                           n8240);
   U10303 : INV_X1 port map( A => ADD_RD1(0), ZN => n6749);
   U10304 : INV_X1 port map( A => ADD_RD2(0), ZN => n6753);
   U10305 : INV_X1 port map( A => ADD_RD1(2), ZN => n6747);
   U10306 : INV_X1 port map( A => ADD_RD2(2), ZN => n6751);
   U10307 : INV_X1 port map( A => ADD_RD1(1), ZN => n6748);
   U10308 : INV_X1 port map( A => ADD_RD2(1), ZN => n6752);
   U10309 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n8274);
   U10310 : AND3_X1 port map( A1 => ENABLE, A2 => n6742, A3 => WR, ZN => n8237)
                           ;
   U10311 : INV_X1 port map( A => ADD_WR(4), ZN => n6742);
   U10312 : INV_X1 port map( A => ADD_WR(3), ZN => n6743);
   U10313 : INV_X1 port map( A => ADD_WR(2), ZN => n6744);
   U10314 : NOR2_X1 port map( A1 => RESET, A2 => n9684, ZN => n8323);
   U10315 : NOR2_X1 port map( A1 => RESET, A2 => n10078, ZN => n7655);
   U10316 : INV_X1 port map( A => RESET, ZN => n6741);
   U10317 : INV_X1 port map( A => DATAIN(0), ZN => n6785);
   U10318 : INV_X1 port map( A => DATAIN(1), ZN => n6784);
   U10319 : INV_X1 port map( A => DATAIN(2), ZN => n6783);
   U10320 : INV_X1 port map( A => DATAIN(3), ZN => n6782);
   U10321 : INV_X1 port map( A => DATAIN(4), ZN => n6781);
   U10322 : INV_X1 port map( A => DATAIN(5), ZN => n6780);
   U10323 : INV_X1 port map( A => DATAIN(6), ZN => n6779);
   U10324 : INV_X1 port map( A => DATAIN(7), ZN => n6778);
   U10325 : INV_X1 port map( A => DATAIN(8), ZN => n6777);
   U10326 : INV_X1 port map( A => DATAIN(9), ZN => n6776);
   U10327 : INV_X1 port map( A => DATAIN(10), ZN => n6775);
   U10328 : INV_X1 port map( A => DATAIN(11), ZN => n6774);
   U10329 : INV_X1 port map( A => DATAIN(12), ZN => n6773);
   U10330 : INV_X1 port map( A => DATAIN(13), ZN => n6772);
   U10331 : INV_X1 port map( A => DATAIN(14), ZN => n6771);
   U10332 : INV_X1 port map( A => DATAIN(15), ZN => n6770);
   U10333 : INV_X1 port map( A => DATAIN(16), ZN => n6769);
   U10334 : INV_X1 port map( A => DATAIN(17), ZN => n6768);
   U10335 : INV_X1 port map( A => DATAIN(18), ZN => n6767);
   U10336 : INV_X1 port map( A => DATAIN(19), ZN => n6766);
   U10337 : INV_X1 port map( A => DATAIN(20), ZN => n6765);
   U10338 : INV_X1 port map( A => DATAIN(21), ZN => n6764);
   U10339 : INV_X1 port map( A => DATAIN(22), ZN => n6763);
   U10340 : INV_X1 port map( A => DATAIN(23), ZN => n6762);
   U10341 : INV_X1 port map( A => DATAIN(24), ZN => n6761);
   U10342 : INV_X1 port map( A => DATAIN(25), ZN => n6760);
   U10343 : INV_X1 port map( A => DATAIN(26), ZN => n6759);
   U10344 : INV_X1 port map( A => DATAIN(27), ZN => n6758);
   U10345 : INV_X1 port map( A => DATAIN(28), ZN => n6757);
   U10346 : INV_X1 port map( A => DATAIN(29), ZN => n6756);
   U10347 : INV_X1 port map( A => DATAIN(30), ZN => n6755);
   U10348 : INV_X1 port map( A => DATAIN(31), ZN => n6754);
   U10349 : INV_X1 port map( A => ADD_RD1(3), ZN => n6746);
   U10350 : INV_X1 port map( A => ADD_RD2(3), ZN => n6750);
   U10351 : INV_X1 port map( A => ADD_WR(0), ZN => n6745);

end SYN_BEHAVIORAL;
