package rf_pkg;
    import uvm_pkg::*;
    import rf_parameters::*;
    `include "uvm_macros.svh"
    `include "data_packet.sv"
    `include "rf_driver.sv"
    `include "rf_monitor.sv"
    `include "rf_sequencer.sv"
    `include "rf_agent.sv"
    `include "rf_scoreboard.sv"
    `include "rf_coverage.sv"
    `include "rf_env.sv"
    `include "dut_env.sv"
    `include "rf_sequences.sv"
    `include "tests.sv"

endpackage