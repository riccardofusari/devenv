class coverage extends uvm_component;
`uvm_component_utils(coverage);

    function new();
        
    endfunction //new()
endclass //coverage extends uvm_component